logic [15:0] rnd_biases [41:0] = { 16'b0011001110110100,	//6.462664
								   16'b0010111110111000,	//5.964799 
								   16'b0001011010011111,	//2.827580 
								   16'b0000001011010001,	//0.352154 
								   16'b1111100110010011,	//-0.803025 
								   16'b0011011010000001,	//6.813164 
								   16'b1110010000001000,	//-3.495889 
								   16'b1110011010000101,	//-3.184913 
								   16'b1110001001010100,	//-3.709082 
								   16'b1111101111111111,	//-0.500447 
								   16'b0000011011100101,	//0.861658 
								   16'b1111111000010100,	//-0.240202 
								   16'b0010000100000010,	//4.126099 
								   16'b0011001011001010,	//6.348553 
								   16'b0000111011100101,	//1.861595 
								   16'b0001101010000100,	//3.314213 
								   16'b0000100100001110,	//1.132060 
								   16'b0000010010010101,	//0.572859 
								   16'b0000000100100011,	//0.142093 
								   16'b1111000101011110,	//-1.829067 
								   16'b1110000011000011,	//-3.904630 
								   16'b1111110011110111,	//-0.379339 
								   16'b0010010000100000,	//4.515650 
								   16'b0001101010000111,	//3.315736 
								   16'b1111101011001010,	//-0.651412 
								   16'b0000011000100101,	//0.767910 
								   16'b0001000001111000,	//2.058438 
								   16'b0000100001101010,	//1.051864 
								   16'b0000011110111101,	//0.967526 
								   16'b0001011010110100,	//2.837687 
								   16'b0000001001110010,	//0.305544 
								   16'b1110101000100101,	//-2.731722 
								   16'b1111000101000001,	//-1.843131 
								   16'b1110100110000100,	//-2.810365 
								   16'b1101111001010101,	//-4.208594 
								   16'b1110100000000011,	//-2.998569 
								   16'b1100110001111000,	//-6.441420 
								   16'b1101001010100001,	//-5.671507 
								   16'b1110010111100011,	//-3.264375 
								   16'b0001000101001100,	//2.162152 
								   16'b1101110100010011,	//-4.365597 
								   16'b1101100101001010};	//-4.838783 

logic [15:0] rnd_inputs [783:0] = {16'b0000100011110111,	//1.120702
								   16'b1111101011001101,	//-0.649665 
								   16'b0000001101110100,	//0.431464 
								   16'b0000011110111000,	//0.965016 
								   16'b1111001101011011,	//-1.580747 
								   16'b1111010000011000,	//-1.488446 
								   16'b0000000110010110,	//0.198160 
								   16'b1111111110000111,	//-0.059082 
								   16'b0000110001111111,	//1.561903 
								   16'b0000100110010001,	//1.195841 
								   16'b0000011110000000,	//0.937364 
								   16'b1111000110100101,	//-1.794672 
								   16'b1111001001010101,	//-1.708459 
								   16'b1111001011010101,	//-1.645890 
								   16'b0000100110001100,	//1.193403 
								   16'b0000111000101101,	//1.772033 
								   16'b0000010111100001,	//0.734862 
								   16'b1111010000111010,	//-1.471668 
								   16'b0000011100100001,	//0.890898 
								   16'b1111001110001000,	//-1.558586 
								   16'b1111001111000011,	//-1.530029 
								   16'b0000010010000001,	//0.562872 
								   16'b1111101010000110,	//-0.684743 
								   16'b0000010011101100,	//0.615248 
								   16'b0000011111111001,	//0.996526 
								   16'b0000001010101001,	//0.332743 
								   16'b0000011110101110,	//0.960129 
								   16'b1111011110000100,	//-1.060692 
								   16'b0000011110000101,	//0.939830 
								   16'b0000111100001111,	//1.882394 
								   16'b0000101110111110,	//1.467721 
								   16'b1111001011000010,	//-1.655062 
								   16'b1111101110111010,	//-0.534254 
								   16'b1111101111010000,	//-0.523205 
								   16'b0000010111101100,	//0.740114 
								   16'b0000001100100010,	//0.391767 
								   16'b0000100101000010,	//1.157456 
								   16'b1111101111000100,	//-0.529388 
								   16'b1111011010011000,	//-1.175889 
								   16'b1111001011000110,	//-1.653334 
								   16'b0000100010110100,	//1.087736 
								   16'b1111011010010101,	//-1.177302 
								   16'b1111110001101101,	//-0.446913 
								   16'b0000000110101000,	//0.207114 
								   16'b1111011101010100,	//-1.084187 
								   16'b0000010010001011,	//0.567762 
								   16'b1111111110000001,	//-0.062079 
								   16'b1111010011011100,	//-1.392618 
								   16'b0000100100000110,	//1.127728 
								   16'b1111001100111000,	//-1.597575 
								   16'b1111100101101001,	//-0.823735 
								   16'b1111011110011001,	//-1.050508 
								   16'b0000000011111101,	//0.123489 
								   16'b1111001011101110,	//-1.634005 
								   16'b1111110011111000,	//-0.378738 
								   16'b1111001101011011,	//-1.580615 
								   16'b1111001110011000,	//-1.550864 
								   16'b0000100100011010,	//1.137712 
								   16'b1111100101010101,	//-0.833719 
								   16'b0000001101010000,	//0.414134 
								   16'b0000111011011101,	//1.857691 
								   16'b1111110111010111,	//-0.270060 
								   16'b0000011000111011,	//0.779009 
								   16'b0000100001000010,	//1.032397 
								   16'b1111110111011000,	//-0.269431 
								   16'b0000010011111010,	//0.621992 
								   16'b1111001110000011,	//-1.560980 
								   16'b0000110111100001,	//1.735039 
								   16'b1111011000000000,	//-1.250157 
								   16'b1111100010000101,	//-0.935285 
								   16'b0000100110001000,	//1.191321 
								   16'b1111111110011010,	//-0.049585 
								   16'b0000100010011011,	//1.075833 
								   16'b1111110010101100,	//-0.415973 
								   16'b1111100010111100,	//-0.908245 
								   16'b1111000100110001,	//-1.851061 
								   16'b0000010110001100,	//0.693180 
								   16'b1111110110111111,	//-0.281742 
								   16'b1111111001110101,	//-0.193043 
								   16'b0000001110000100,	//0.439429 
								   16'b1111000111100111,	//-1.762387 
								   16'b1111101000011011,	//-0.736754 
								   16'b0000100010111010,	//1.090889 
								   16'b0000011001001001,	//0.785732 
								   16'b1111010000000011,	//-1.498671 
								   16'b1111010000101010,	//-1.479394 
								   16'b1111001011110101,	//-1.630591 
								   16'b1111000001000000,	//-1.968719 
								   16'b1111110110001010,	//-0.307562 
								   16'b0000010011111010,	//0.622293 
								   16'b0000011100100010,	//0.891690 
								   16'b0000000100000000,	//0.124837 
								   16'b1111001101111011,	//-1.564728 
								   16'b0000010000110111,	//0.527065 
								   16'b1111010000001100,	//-1.494001 
								   16'b1111010001001100,	//-1.462787 
								   16'b1111001100101000,	//-1.605624 
								   16'b1111010010001011,	//-1.431891 
								   16'b1111010101100010,	//-1.326995 
								   16'b1111011001001000,	//-1.215004 
								   16'b1111101000101001,	//-0.730081 
								   16'b1111101000100000,	//-0.734284 
								   16'b1111011011110110,	//-1.129747 
								   16'b1111100000001001,	//-0.995833 
								   16'b0000110010010011,	//1.571690 
								   16'b0000011010000001,	//0.812893 
								   16'b0000000111001001,	//0.222952 
								   16'b1111010111100111,	//-1.262265 
								   16'b1111011011001001,	//-1.151877 
								   16'b1111001001111010,	//-1.690613 
								   16'b0000110100111110,	//1.655202 
								   16'b0000011010011101,	//0.826861 
								   16'b0000000111011001,	//0.231156 
								   16'b1111101000001000,	//-0.746284 
								   16'b1111010101010010,	//-1.335186 
								   16'b0000001111101011,	//0.489989 
								   16'b0000111110011101,	//1.951739 
								   16'b1111010101110100,	//-1.318272 
								   16'b1111100001000000,	//-0.968831 
								   16'b1111110010110011,	//-0.412803 
								   16'b1111001001011110,	//-1.704021 
								   16'b0000010111100100,	//0.736384 
								   16'b1111110011100000,	//-0.390447 
								   16'b0000111101110011,	//1.931341 
								   16'b1111110011011111,	//-0.391264 
								   16'b0000001111011101,	//0.482688 
								   16'b1111010011110001,	//-1.382521 
								   16'b1111110000110100,	//-0.474619 
								   16'b1111010100101000,	//-1.355464 
								   16'b0000100001000010,	//1.032450 
								   16'b0000101111100000,	//1.484444 
								   16'b1111101100111010,	//-0.596893 
								   16'b0000010111110000,	//0.742143 
								   16'b1111100101101010,	//-0.823405 
								   16'b0000000011111011,	//0.122517 
								   16'b0000101010100011,	//1.329694 
								   16'b0000001100011111,	//0.389961 
								   16'b1111101010111011,	//-0.658755 
								   16'b1111100110010011,	//-0.803100 
								   16'b1111111001111100,	//-0.189630 
								   16'b1111110110000110,	//-0.309417 
								   16'b1111101110000010,	//-0.561575 
								   16'b0000000111011110,	//0.233277 
								   16'b0000011111000011,	//0.970181 
								   16'b1111110110010100,	//-0.302661 
								   16'b1111110110111101,	//-0.282577 
								   16'b1111001111111111,	//-1.500509 
								   16'b1111000011001000,	//-1.902264 
								   16'b1111100101001001,	//-0.839259 
								   16'b1111101000101001,	//-0.729918 
								   16'b0000010011101011,	//0.614761 
								   16'b0000111010011111,	//1.827744 
								   16'b0000110111110010,	//1.742923 
								   16'b1111111010100111,	//-0.168455 
								   16'b1111011110110010,	//-1.038086 
								   16'b0000100001110010,	//1.055592 
								   16'b0000100001001100,	//1.037310 
								   16'b0000011110110011,	//0.962592 
								   16'b0000011111001100,	//0.974753 
								   16'b1111001101100100,	//-1.576318 
								   16'b0000010111001111,	//0.726242 
								   16'b1111111011010011,	//-0.146958 
								   16'b1111011011001010,	//-1.151347 
								   16'b1111001100100111,	//-1.605925 
								   16'b0000101001011011,	//1.294298 
								   16'b1111010110011010,	//-1.299961 
								   16'b1111010100111100,	//-1.345720 
								   16'b0000010101010000,	//0.663949 
								   16'b0000110010011111,	//1.577558 
								   16'b0000000010001000,	//0.066233 
								   16'b0000011001111101,	//0.810809 
								   16'b1111010011101010,	//-1.385638 
								   16'b0000111010000011,	//1.813828 
								   16'b0000000101001111,	//0.163536 
								   16'b0000010111000000,	//0.718936 
								   16'b1111000100101100,	//-1.853748 
								   16'b0000100111100101,	//1.236815 
								   16'b0000011111110101,	//0.994475 
								   16'b1111001111011001,	//-1.519252 
								   16'b0000000011001101,	//0.100181 
								   16'b1111101001101101,	//-0.696665 
								   16'b0000000101111101,	//0.185798 
								   16'b1111110011000100,	//-0.404477 
								   16'b1111110101001000,	//-0.339626 
								   16'b1111010111001001,	//-1.277049 
								   16'b1111100000101100,	//-0.978453 
								   16'b1111000010101000,	//-1.917857 
								   16'b0000110110001111,	//1.694702 
								   16'b0000010011101011,	//0.614800 
								   16'b0000110111011000,	//1.730454 
								   16'b1111010100111011,	//-1.345951 
								   16'b0000110101111010,	//1.684389 
								   16'b0000100101101110,	//1.178632 
								   16'b0000001001111010,	//0.309577 
								   16'b1111111000010101,	//-0.239858 
								   16'b1111100000111110,	//-0.969545 
								   16'b0000100000010000,	//1.007786 
								   16'b1111011101010001,	//-1.085322 
								   16'b1111001000001110,	//-1.743252 
								   16'b0000100010001110,	//1.069318 
								   16'b0000010101111010,	//0.684809 
								   16'b0000011011100011,	//0.860850 
								   16'b0000010010001100,	//0.568243 
								   16'b1111110101101001,	//-0.323807 
								   16'b1111110010000001,	//-0.436952 
								   16'b0000101000011110,	//1.264560 
								   16'b1111101000101000,	//-0.730289 
								   16'b0000101000010001,	//1.258159 
								   16'b0000100101000000,	//1.156294 
								   16'b0000101101000110,	//1.409056 
								   16'b0000000000101110,	//0.022546 
								   16'b0000010001010111,	//0.542646 
								   16'b0000111001101110,	//1.803578 
								   16'b1111111000110101,	//-0.224143 
								   16'b1111000111101100,	//-1.759925 
								   16'b0000101110111100,	//1.467000 
								   16'b0000010000110011,	//0.524755 
								   16'b1111101101011101,	//-0.579705 
								   16'b0000111111100111,	//1.988013 
								   16'b1111011100101100,	//-1.103314 
								   16'b0000010011100001,	//0.609804 
								   16'b0000001101011100,	//0.419963 
								   16'b1111110001100100,	//-0.451018 
								   16'b1111010010001101,	//-1.431251 
								   16'b1111000011001110,	//-1.899460 
								   16'b1111110101111010,	//-0.315551 
								   16'b1111010111100100,	//-1.263599 
								   16'b0000011100111010,	//0.903101 
								   16'b1111101111011010,	//-0.518549 
								   16'b0000101011101110,	//1.366240 
								   16'b0000011101111111,	//0.936919 
								   16'b0000001001000110,	//0.284103 
								   16'b1111010110101001,	//-1.292580 
								   16'b0000111010100011,	//1.829536 
								   16'b1111100001111110,	//-0.938712 
								   16'b0000110110010110,	//1.698324 
								   16'b1111011100101001,	//-1.104918 
								   16'b1111101111110100,	//-0.505745 
								   16'b1111001011001101,	//-1.649999 
								   16'b0000010001111100,	//0.560466 
								   16'b1111010111001000,	//-1.277532 
								   16'b1111000101110001,	//-1.819796 
								   16'b0000011100100100,	//0.892694 
								   16'b1111101100011110,	//-0.610249 
								   16'b0000010100100100,	//0.642467 
								   16'b1111110001001001,	//-0.464526 
								   16'b0000010000010011,	//0.509386 
								   16'b1111000010110001,	//-1.913401 
								   16'b0000110100100011,	//1.642280 
								   16'b0000100110011110,	//1.202235 
								   16'b0000011111011110,	//0.983390 
								   16'b0000101000000101,	//1.252451 
								   16'b1111110001000100,	//-0.466775 
								   16'b0000001111000001,	//0.469117 
								   16'b0000001001101010,	//0.301979 
								   16'b0000000011110110,	//0.120207 
								   16'b1111100011001101,	//-0.899721 
								   16'b1111011111110101,	//-1.005484 
								   16'b1111111001110100,	//-0.193445 
								   16'b1111011101001001,	//-1.089149 
								   16'b0000100110111110,	//1.217798 
								   16'b0000111110001110,	//1.944417 
								   16'b1111000011110110,	//-1.880032 
								   16'b0000000100100100,	//0.142657 
								   16'b1111001011001001,	//-1.651691 
								   16'b0000100110101011,	//1.208366 
								   16'b0000111110100111,	//1.956580 
								   16'b1111001000100100,	//-1.732215 
								   16'b0000111000010000,	//1.757593 
								   16'b1111000010010101,	//-1.927290 
								   16'b0000010111100010,	//0.735354 
								   16'b0000100100010100,	//1.134946 
								   16'b0000000100011000,	//0.136550 
								   16'b0000110001010101,	//1.541438 
								   16'b0000110011000101,	//1.596020 
								   16'b0000010000001000,	//0.503751 
								   16'b1111010001101001,	//-1.448524 
								   16'b1111011011111000,	//-1.128794 
								   16'b1111010111010100,	//-1.271436 
								   16'b1111000101010111,	//-1.832721 
								   16'b1111001101101100,	//-1.572233 
								   16'b0000001110111010,	//0.465774 
								   16'b0000111000010010,	//1.758644 
								   16'b1111101101011000,	//-0.582177 
								   16'b1111110100100100,	//-0.357484 
								   16'b0000111110000000,	//1.937398 
								   16'b0000111001000010,	//1.782317 
								   16'b0000010110100111,	//0.706579 
								   16'b0000111110100000,	//1.953209 
								   16'b0000100010001010,	//1.067326 
								   16'b1111101011000110,	//-0.653203 
								   16'b0000010100110010,	//0.649527 
								   16'b1111011111010000,	//-1.023339 
								   16'b1111100101110101,	//-0.817971 
								   16'b0000010111000100,	//0.720713 
								   16'b0000000011100100,	//0.111387 
								   16'b1111110100101100,	//-0.353626 
								   16'b0000001101001001,	//0.410553 
								   16'b0000100000000100,	//1.002080 
								   16'b0000001010101100,	//0.334133 
								   16'b0000000110101000,	//0.207170 
								   16'b0000001010101101,	//0.334282 
								   16'b0000000001100001,	//0.047280 
								   16'b1111001010100101,	//-1.669629 
								   16'b0000011100000111,	//0.878281 
								   16'b0000111111100001,	//1.984624 
								   16'b1111101101011000,	//-0.581863 
								   16'b0000111100010101,	//1.885035 
								   16'b1111101100010110,	//-0.614205 
								   16'b0000110001011111,	//1.546175 
								   16'b1111111010001101,	//-0.181221 
								   16'b1111110100111011,	//-0.346291 
								   16'b1111011011111000,	//-1.129072 
								   16'b1111010000000101,	//-1.497382 
								   16'b1111100111100011,	//-0.764342 
								   16'b0000011100111100,	//0.904418 
								   16'b0000100100001101,	//1.131488 
								   16'b0000011000110100,	//0.775150 
								   16'b1111000001010000,	//-1.960791 
								   16'b0000101011111100,	//1.372853 
								   16'b0000110110000100,	//1.689328 
								   16'b0000100010101100,	//1.083817 
								   16'b1111000101011101,	//-1.829361 
								   16'b1111110000011010,	//-0.487255 
								   16'b0000011010001010,	//0.817358 
								   16'b0000011101011000,	//0.918052 
								   16'b1111011100101101,	//-1.102892 
								   16'b1111100010011100,	//-0.923781 
								   16'b0000010110001001,	//0.692125 
								   16'b1111111101001000,	//-0.090031 
								   16'b0000001111110101,	//0.494866 
								   16'b1111011110010001,	//-1.054220 
								   16'b1111010110101011,	//-1.291505 
								   16'b0000101010001100,	//1.318574 
								   16'b0000100010001011,	//1.067687 
								   16'b0000110111100111,	//1.737913 
								   16'b1111001101110100,	//-1.568444 
								   16'b1111010111010101,	//-1.271090 
								   16'b1111001100101100,	//-1.603619 
								   16'b1111111110101100,	//-0.040945 
								   16'b1111011000101111,	//-1.227019 
								   16'b0000110010101011,	//1.583566 
								   16'b1111001100101100,	//-1.603641 
								   16'b1111000101101010,	//-1.823338 
								   16'b0000000111010101,	//0.229181 
								   16'b0000100010111000,	//1.089980 
								   16'b1111100111111011,	//-0.752240 
								   16'b1111010110111010,	//-1.284070 
								   16'b1111101011011001,	//-0.644177 
								   16'b1111011010111010,	//-1.159417 
								   16'b0000000001010011,	//0.040610 
								   16'b0000110100000001,	//1.625457 
								   16'b0000010000100000,	//0.515696 
								   16'b1111001101000000,	//-1.593864 
								   16'b1111110010000010,	//-0.436581 
								   16'b1111000110111111,	//-1.781534 
								   16'b0000000000001011,	//0.005132 
								   16'b1111110111010001,	//-0.273115 
								   16'b0000111111101100,	//1.990241 
								   16'b0000100111111001,	//1.246410 
								   16'b1111111110001010,	//-0.057393 
								   16'b0000110010011111,	//1.577791 
								   16'b1111010001100111,	//-1.449814 
								   16'b1111110001111011,	//-0.439980 
								   16'b0000110110101101,	//1.709425 
								   16'b0000110101011100,	//1.669975 
								   16'b0000011011010110,	//0.854296 
								   16'b0000001111001001,	//0.473350 
								   16'b1111101011111100,	//-0.626848 
								   16'b0000110111110100,	//1.744109 
								   16'b1111001111111110,	//-1.500904 
								   16'b0000011101100001,	//0.922341 
								   16'b0000010010110000,	//0.585910 
								   16'b0000101010101001,	//1.332608 
								   16'b1111110010111111,	//-0.406871 
								   16'b0000011111111111,	//0.999289 
								   16'b0000101010111010,	//1.340882 
								   16'b1111101001010010,	//-0.710158 
								   16'b0000000110101100,	//0.209046 
								   16'b0000111101010101,	//1.916517 
								   16'b0000000110010100,	//0.197234 
								   16'b1111101010010011,	//-0.678306 
								   16'b0000001111010011,	//0.477886 
								   16'b1111101110001010,	//-0.557454 
								   16'b0000100000110101,	//1.026038 
								   16'b1111110100111111,	//-0.344397 
								   16'b1111111111000001,	//-0.030620 
								   16'b0000011000111011,	//0.778973 
								   16'b0000111100100001,	//1.890936 
								   16'b1111101001111101,	//-0.688980 
								   16'b0000101011001111,	//1.351213 
								   16'b0000011110100110,	//0.956289 
								   16'b0000111010001001,	//1.816698 
								   16'b1111000100000110,	//-1.872309 
								   16'b1111101101101011,	//-0.572524 
								   16'b0000010100110100,	//0.650615 
								   16'b1111100100000010,	//-0.873994 
								   16'b1111011101011111,	//-1.078468 
								   16'b0000011011000010,	//0.844514 
								   16'b0000001111111101,	//0.498292 
								   16'b0000001011100110,	//0.362435 
								   16'b0000010100100010,	//0.641752 
								   16'b1111000110000110,	//-1.809781 
								   16'b1111101100101001,	//-0.604861 
								   16'b1111111001110001,	//-0.194638 
								   16'b1111011110110101,	//-1.036380 
								   16'b0000011011100010,	//0.860180 
								   16'b0000101101100110,	//1.424729 
								   16'b1111100100000010,	//-0.873969 
								   16'b0000011101100101,	//0.924203 
								   16'b1111010001101001,	//-1.448948 
								   16'b0000101011000110,	//1.346891 
								   16'b1111010001101111,	//-1.445593 
								   16'b0000001011010011,	//0.352838 
								   16'b1111101110111000,	//-0.535373 
								   16'b0000100111010001,	//1.227038 
								   16'b0000000000011111,	//0.015123 
								   16'b1111111110101011,	//-0.041623 
								   16'b0000110000010001,	//1.508195 
								   16'b1111101101001101,	//-0.587433 
								   16'b1111111001100010,	//-0.202226 
								   16'b0000111011010101,	//1.854121 
								   16'b1111000101011011,	//-1.830809 
								   16'b0000111100100010,	//1.891833 
								   16'b1111011000001110,	//-1.243173 
								   16'b0000010101011001,	//0.668481 
								   16'b0000001011000100,	//0.345758 
								   16'b0000010110011011,	//0.700450 
								   16'b1111101110001101,	//-0.555912 
								   16'b0000001111011001,	//0.481114 
								   16'b0000100111110101,	//1.244604 
								   16'b1111000010011110,	//-1.922970 
								   16'b1111001010101111,	//-1.664506 
								   16'b0000111100110010,	//1.899207 
								   16'b0000010011011000,	//0.605398 
								   16'b1111011101100110,	//-1.075049 
								   16'b1111110011101001,	//-0.386035 
								   16'b1111001111101000,	//-1.511918 
								   16'b1111100010010111,	//-0.926245 
								   16'b1111100001000000,	//-0.968615 
								   16'b1111101010011101,	//-0.673339 
								   16'b1111010011011111,	//-1.391064 
								   16'b1111101100100011,	//-0.607969 
								   16'b1111001111100101,	//-1.513366 
								   16'b0000110001001011,	//1.536612 
								   16'b1111001100000100,	//-1.622886 
								   16'b0000110111000011,	//1.720163 
								   16'b1111110011000101,	//-0.403920 
								   16'b1111000110000100,	//-1.810394 
								   16'b1111101011110101,	//-0.630506 
								   16'b0000011110001101,	//0.943865 
								   16'b0000100101101110,	//1.178729 
								   16'b0000000101110000,	//0.179624 
								   16'b0000010111110110,	//0.744894 
								   16'b0000110010011001,	//1.574531 
								   16'b1111000111000001,	//-1.780833 
								   16'b1111100110111000,	//-0.785354 
								   16'b1111000101111010,	//-1.815234 
								   16'b1111011001000001,	//-1.218093 
								   16'b0000011100001100,	//0.880663 
								   16'b0000011100011001,	//0.887013 
								   16'b0000110000010111,	//1.511196 
								   16'b0000001010100011,	//0.329732 
								   16'b1111001001000011,	//-1.717263 
								   16'b0000110110000111,	//1.690978 
								   16'b0000100110011101,	//1.201488 
								   16'b1111100100100110,	//-0.856213 
								   16'b0000000101100110,	//0.174653 
								   16'b0000111110000011,	//1.939105 
								   16'b0000011011100111,	//0.862712 
								   16'b0000101011011001,	//1.355878 
								   16'b1111110111011101,	//-0.266958 
								   16'b1111111100001111,	//-0.117501 
								   16'b0000000111110001,	//0.242854 
								   16'b1111100010011100,	//-0.923634 
								   16'b0000011111111000,	//0.996074 
								   16'b0000000000100000,	//0.015551 
								   16'b0000010010110011,	//0.587239 
								   16'b1111100111011001,	//-0.769018 
								   16'b1111010001110000,	//-1.445101 
								   16'b1111111100111000,	//-0.097708 
								   16'b1111101110011001,	//-0.550163 
								   16'b0000100100111000,	//1.152454 
								   16'b0000100011111000,	//1.121183 
								   16'b0000010101100100,	//0.674049 
								   16'b1111010001000110,	//-1.465985 
								   16'b1111000010110001,	//-1.913776 
								   16'b0000000111101010,	//0.239363 
								   16'b1111100110100000,	//-0.796724 
								   16'b0000111000010000,	//1.757639 
								   16'b0000111101100100,	//1.923615 
								   16'b1111100100101100,	//-0.853518 
								   16'b0000100110100000,	//1.203281 
								   16'b0000110010101101,	//1.584445 
								   16'b0000001100011111,	//0.390106 
								   16'b0000110001001010,	//1.536067 
								   16'b0000111000110011,	//1.774926 
								   16'b0000000110010011,	//0.196632 
								   16'b0000011101001111,	//0.913547 
								   16'b0000001001110101,	//0.307033 
								   16'b1111000011010100,	//-1.896570 
								   16'b1111111001001010,	//-0.213876 
								   16'b0000010010101111,	//0.585208 
								   16'b0000000010101110,	//0.084812 
								   16'b1111101111101010,	//-0.510749 
								   16'b0000110111111101,	//1.748539 
								   16'b0000101010001100,	//1.318131 
								   16'b0000101100101100,	//1.396342 
								   16'b1111101111101100,	//-0.509863 
								   16'b0000001011111011,	//0.372738 
								   16'b0000101111101100,	//1.490210 
								   16'b0000110111011111,	//1.734006 
								   16'b0000010101100100,	//0.673857 
								   16'b1111011010011110,	//-1.172894 
								   16'b0000010011101100,	//0.615402 
								   16'b1111001001001110,	//-1.711794 
								   16'b1111110100000100,	//-0.373092 
								   16'b0000010101011000,	//0.667726 
								   16'b0000110111100001,	//1.734903 
								   16'b0000100111110011,	//1.243800 
								   16'b1111111110000001,	//-0.061807 
								   16'b0000100000110111,	//1.026997 
								   16'b1111110101011000,	//-0.331810 
								   16'b0000111100011001,	//1.887144 
								   16'b0000111110011101,	//1.951899 
								   16'b0000101110100111,	//1.456590 
								   16'b1111110001110010,	//-0.444465 
								   16'b1111111010001101,	//-0.181033 
								   16'b1111011111100101,	//-1.013251 
								   16'b0000100100011010,	//1.137692 
								   16'b0000110001000000,	//1.531350 
								   16'b0000110100111101,	//1.654847 
								   16'b0000000111011101,	//0.233140 
								   16'b0000001100101010,	//0.395472 
								   16'b1111010011000100,	//-1.404493 
								   16'b0000110011001010,	//1.598854 
								   16'b1111111001101010,	//-0.198426 
								   16'b1111011010010101,	//-1.177311 
								   16'b0000110011001010,	//1.598604 
								   16'b0000100001100111,	//1.050342 
								   16'b0000110000111101,	//1.529945 
								   16'b1111100100011110,	//-0.860199 
								   16'b0000010110001011,	//0.692904 
								   16'b0000010101000010,	//0.657120 
								   16'b1111001111101110,	//-1.508740 
								   16'b1111110100001001,	//-0.370726 
								   16'b1111100011001111,	//-0.898852 
								   16'b0000011011101111,	//0.866679 
								   16'b1111100100010001,	//-0.866462 
								   16'b0000110010101110,	//1.584795 
								   16'b0000101001110011,	//1.306316 
								   16'b1111110001111011,	//-0.439894 
								   16'b1111111111101111,	//-0.008388 
								   16'b0000011000111100,	//0.779221 
								   16'b0000101010110011,	//1.337476 
								   16'b0000001110000010,	//0.438519 
								   16'b0000001001100100,	//0.298949 
								   16'b1111101001101111,	//-0.695831 
								   16'b1111111010011011,	//-0.174302 
								   16'b0000011011010111,	//0.855182 
								   16'b0000110001001101,	//1.537620 
								   16'b0000011100010001,	//0.883423 
								   16'b1111000010011000,	//-1.925549 
								   16'b0000010110011000,	//0.699106 
								   16'b1111111000001000,	//-0.245965 
								   16'b1111111000000011,	//-0.248719 
								   16'b1111001110111111,	//-1.531853 
								   16'b0000101000010010,	//1.258727 
								   16'b1111101001100101,	//-0.700578 
								   16'b1111011111100001,	//-1.015088 
								   16'b1111101011111000,	//-0.629147 
								   16'b1111110000000110,	//-0.497231 
								   16'b0000000101111101,	//0.186215 
								   16'b0000000111111011,	//0.247681 
								   16'b1111110010101011,	//-0.416711 
								   16'b1111110010111101,	//-0.407476 
								   16'b0000000001111110,	//0.061469 
								   16'b0000010100001010,	//0.630122 
								   16'b0000111001101110,	//1.803661 
								   16'b0000011100011101,	//0.889394 
								   16'b1111110011001101,	//-0.399681 
								   16'b0000101010011111,	//1.327485 
								   16'b1111010001001100,	//-1.462647 
								   16'b1111000111101111,	//-1.758133 
								   16'b1111001010110010,	//-1.663012 
								   16'b1111010100111111,	//-1.344407 
								   16'b1111101001100000,	//-0.703120 
								   16'b1111100110101000,	//-0.793093 
								   16'b1111000001100000,	//-1.953276 
								   16'b0000000101000111,	//0.159620 
								   16'b1111001100001101,	//-1.618509 
								   16'b1111010010110000,	//-1.413941 
								   16'b0000010000110010,	//0.524565 
								   16'b0000101110000000,	//1.437282 
								   16'b0000111100101101,	//1.896887 
								   16'b0000001001000100,	//0.283354 
								   16'b0000111111100110,	//1.987401 
								   16'b0000000110110111,	//0.214166 
								   16'b0000000001111111,	//0.061834 
								   16'b1111101010010101,	//-0.677272 
								   16'b1111110111000011,	//-0.279993 
								   16'b1111111110111101,	//-0.032775 
								   16'b1111001001000110,	//-1.715852 
								   16'b0000110001101000,	//1.550957 
								   16'b1111001000010001,	//-1.741466 
								   16'b1111110111110101,	//-0.255260 
								   16'b0000101001110100,	//1.306518 
								   16'b1111110010100000,	//-0.421861 
								   16'b0000001110100010,	//0.453900 
								   16'b0000101000110010,	//1.274563 
								   16'b0000110001011100,	//1.544940 
								   16'b0000110111001100,	//1.724447 
								   16'b1111011000011011,	//-1.236861 
								   16'b1111100001000110,	//-0.965671 
								   16'b0000110010111011,	//1.591463 
								   16'b0000001011111101,	//0.373447 
								   16'b0000000000011111,	//0.015360 
								   16'b0000001110011100,	//0.451238 
								   16'b0000101000111001,	//1.277689 
								   16'b0000000100000101,	//0.127557 
								   16'b1111011001110111,	//-1.191700 
								   16'b1111111010000110,	//-0.184426 
								   16'b1111110110110001,	//-0.288356 
								   16'b0000111011101010,	//1.864211 
								   16'b0000001111010111,	//0.480220 
								   16'b0000011001000001,	//0.781560 
								   16'b0000011100001100,	//0.880658 
								   16'b1111101100011010,	//-0.612419 
								   16'b0000000010001011,	//0.067962 
								   16'b0000000111010000,	//0.226779 
								   16'b1111010100000010,	//-1.374019 
								   16'b0000000111111100,	//0.248224 
								   16'b0000011000111100,	//0.779213 
								   16'b1111110110100110,	//-0.294178 
								   16'b0000101011000011,	//1.345082 
								   16'b0000011101101000,	//0.925548 
								   16'b1111101110000101,	//-0.559876 
								   16'b1111111010001001,	//-0.183151 
								   16'b1111110001011101,	//-0.454440 
								   16'b0000100011010001,	//1.102219 
								   16'b0000011101111111,	//0.937084 
								   16'b1111110111000101,	//-0.278889 
								   16'b0000011000110011,	//0.775010 
								   16'b0000111000111111,	//1.780854 
								   16'b0000100100011000,	//1.136930 
								   16'b0000011010010100,	//0.822287 
								   16'b1111001110000000,	//-1.562663 
								   16'b1111110001111010,	//-0.440277 
								   16'b0000001011101001,	//0.363619 
								   16'b1111111010110011,	//-0.162480 
								   16'b1111000110011100,	//-1.798640 
								   16'b1111011101010001,	//-1.085250 
								   16'b0000101010110010,	//1.336756 
								   16'b1111000010000000,	//-1.937421 
								   16'b0000101110100100,	//1.454843 
								   16'b1111001010000000,	//-1.687724 
								   16'b0000010101101001,	//0.676170 
								   16'b0000000000000010,	//0.000845 
								   16'b1111011011111010,	//-1.128025 
								   16'b0000001001001011,	//0.286463 
								   16'b1111001111101001,	//-1.511243 
								   16'b0000010101111010,	//0.684665 
								   16'b0000001100110000,	//0.398342 
								   16'b1111000111001011,	//-1.776095 
								   16'b1111000111001110,	//-1.774628 
								   16'b1111010011100001,	//-1.389997 
								   16'b1111000010100001,	//-1.921516 
								   16'b1111110111101101,	//-0.259298 
								   16'b0000101010100010,	//1.328886 
								   16'b0000001111000010,	//0.469561 
								   16'b0000000010100101,	//0.080518 
								   16'b0000101110100101,	//1.455473 
								   16'b1111001100100000,	//-1.609208 
								   16'b0000110100001111,	//1.632209 
								   16'b1111001101110101,	//-1.567933 
								   16'b0000000010001011,	//0.067987 
								   16'b1111010010010101,	//-1.427376 
								   16'b0000000111100110,	//0.237482 
								   16'b1111000000100110,	//-1.981682 
								   16'b0000100010001001,	//1.066728 
								   16'b0000101100101001,	//1.394837 
								   16'b0000110101010111,	//1.667285 
								   16'b0000111110010101,	//1.947873 
								   16'b0000000000101010,	//0.020532 
								   16'b1111100010101111,	//-0.914314 
								   16'b1111001100111001,	//-1.596998 
								   16'b0000000001000000,	//0.031395 
								   16'b0000001010111101,	//0.342437 
								   16'b0000100001101010,	//1.051548 
								   16'b1111001010101000,	//-1.668149 
								   16'b0000010100101100,	//0.646385 
								   16'b0000000010001011,	//0.067916 
								   16'b1111010101111001,	//-1.315808 
								   16'b0000111000001001,	//1.754231 
								   16'b0000001011100101,	//0.361933 
								   16'b1111111000011010,	//-0.237461 
								   16'b0000111000100100,	//1.767676 
								   16'b0000010011111101,	//0.623655 
								   16'b1111111001110110,	//-0.192217 
								   16'b0000101011011111,	//1.358790 
								   16'b0000000100001011,	//0.130494 
								   16'b0000000110111001,	//0.215548 
								   16'b0000010111000011,	//0.720262 
								   16'b1111101111000000,	//-0.531240 
								   16'b1111011110101000,	//-1.042838 
								   16'b0000001010000111,	//0.315694 
								   16'b0000101110111110,	//1.467548 
								   16'b1111110100000100,	//-0.372893 
								   16'b1111001110011011,	//-1.549539 
								   16'b1111111000110100,	//-0.224617 
								   16'b1111100110011011,	//-0.799262 
								   16'b1111110011011000,	//-0.394453 
								   16'b0000101010101011,	//1.333454 
								   16'b1111110011101011,	//-0.385485 
								   16'b1111110001111100,	//-0.439296 
								   16'b1111101110001001,	//-0.558204 
								   16'b1111010001111101,	//-1.438979 
								   16'b1111100001010011,	//-0.959479 
								   16'b1111001011000111,	//-1.652740 
								   16'b1111110110111110,	//-0.282411 
								   16'b1111100000111100,	//-0.970869 
								   16'b1111100110000110,	//-0.809778 
								   16'b1111110110011000,	//-0.300566 
								   16'b1111001111010001,	//-1.523171 
								   16'b1111111111011000,	//-0.019732 
								   16'b0000011010011011,	//0.825629 
								   16'b1111011111001011,	//-1.025707 
								   16'b0000100100011111,	//1.140280 
								   16'b1111001001011111,	//-1.703642 
								   16'b1111110010011011,	//-0.424466 
								   16'b1111000000011100,	//-1.986424 
								   16'b1111011100010000,	//-1.117292 
								   16'b1111000000001011,	//-1.994798 
								   16'b1111011000001110,	//-1.243281 
								   16'b1111010010001111,	//-1.430064 
								   16'b1111100010010100,	//-0.927696 
								   16'b1111010110011001,	//-1.300432 
								   16'b1111010001110000,	//-1.445404 
								   16'b0000001100101010,	//0.395542 
								   16'b0000110011010101,	//1.604232 
								   16'b0000111000001111,	//1.757519 
								   16'b1111011100010100,	//-1.115262 
								   16'b1111111101110010,	//-0.069314 
								   16'b1111110000001000,	//-0.495956 
								   16'b0000000011000011,	//0.095120 
								   16'b1111100001111010,	//-0.940510 
								   16'b1111001000110000,	//-1.726571 
								   16'b1111110111110110,	//-0.254692 
								   16'b1111010110010000,	//-1.304588 
								   16'b1111000011010110,	//-1.895572 
								   16'b0000111010001101,	//1.818713 
								   16'b1111110111000111,	//-0.277614 
								   16'b0000111011000101,	//1.846234 
								   16'b0000100001100110,	//1.049658 
								   16'b1111000000111100,	//-1.970605 
								   16'b0000010111000011,	//0.720155 
								   16'b0000011010010111,	//0.823803 
								   16'b0000010010100101,	//0.580515 
								   16'b0000000110101101,	//0.209239 
								   16'b1111011011111011,	//-1.127565 
								   16'b0000100010110111,	//1.089465 
								   16'b1111011101001100,	//-1.087887 
								   16'b1111101111011110,	//-0.516541 
								   16'b0000110010000010,	//1.563715 
								   16'b0000101101100111,	//1.425508 
								   16'b1111110011100001,	//-0.390266 
								   16'b1111101000101101,	//-0.727924 
								   16'b0000001101111010,	//0.434542 
								   16'b0000110100100000,	//1.640781 
								   16'b0000110100010111,	//1.636393 
								   16'b0000001011101110,	//0.366378 
								   16'b1111101010100100,	//-0.669714 
								   16'b0000101101001100,	//1.412255 
								   16'b1111111000101000,	//-0.230408 
								   16'b0000110011110000,	//1.617422 
								   16'b1111000100010000,	//-1.867282 
								   16'b0000000100001010,	//0.129706 
								   16'b0000011011101110,	//0.865989 
								   16'b1111010110111101,	//-1.282793 
								   16'b1111101011000101,	//-0.653868 
								   16'b1111011000000010,	//-1.249148 
								   16'b1111101001001101,	//-0.712291 
								   16'b1111110011101100,	//-0.384573 
								   16'b0000000110001110};	//0.194265 


logic [15:0] rnd_weights [783:0] = {16'b0000101000010010,	//1.258895 
								   16'b0000110011111100,	//1.623168 
								   16'b1111010000010000,	//-1.492053 
								   16'b0000110100111010,	//1.653503 
								   16'b0000010000111100,	//0.529437 
								   16'b1111001100011111,	//-1.609838 
								   16'b1111100011101001,	//-0.886007 
								   16'b0000000110000000,	//0.187526 
								   16'b0000111010100100,	//1.830027 
								   16'b0000111011100000,	//1.859554 
								   16'b1111010100001011,	//-1.369548 
								   16'b0000111100001111,	//1.882371 
								   16'b0000111010100001,	//1.828668 
								   16'b1111111110001000,	//-0.058497 
								   16'b0000100110011100,	//1.201122 
								   16'b1111010010001010,	//-1.432455 
								   16'b1111110101111111,	//-0.312955 
								   16'b0000110101001110,	//1.662942 
								   16'b0000100101011010,	//1.168829 
								   16'b0000111010110100,	//1.837970 
								   16'b0000010011111100,	//0.622963 
								   16'b1111000100100101,	//-1.857153 
								   16'b0000101100101100,	//1.396517 
								   16'b0000110111100011,	//1.735973 
								   16'b0000010110111000,	//0.714941 
								   16'b0000100000111111,	//1.030961 
								   16'b0000011111001000,	//0.972530 
								   16'b1111110010001101,	//-0.431092 
								   16'b0000010011111010,	//0.621912 
								   16'b1111010101111010,	//-1.315253 
								   16'b0000011010011000,	//0.824184 
								   16'b1111000100000101,	//-1.872669 
								   16'b1111100011011101,	//-0.892308 
								   16'b1111000101111010,	//-1.815314 
								   16'b1111001100011100,	//-1.611473 
								   16'b0000101001011010,	//1.293831 
								   16'b0000011000111100,	//0.779314 
								   16'b1111101000100110,	//-0.731602 
								   16'b0000111001101000,	//1.800888 
								   16'b1111000100011010,	//-1.862216 
								   16'b1111111000001010,	//-0.245023 
								   16'b1111110000110110,	//-0.473766 
								   16'b0000100001111111,	//1.062067 
								   16'b0000100101110010,	//1.180800 
								   16'b1111010111111011,	//-1.252510 
								   16'b1111111110101100,	//-0.040942 
								   16'b1111111001000010,	//-0.217655 
								   16'b0000010010101111,	//0.585252 
								   16'b0000011010110011,	//0.837459 
								   16'b0000100000100110,	//1.018747 
								   16'b1111100011010101,	//-0.895900 
								   16'b0000010111000000,	//0.718811 
								   16'b0000010011110111,	//0.620392 
								   16'b1111010100110100,	//-1.349553 
								   16'b1111001111001111,	//-1.524009 
								   16'b1111111111110011,	//-0.006544 
								   16'b0000111010110110,	//1.838976 
								   16'b1111101011100100,	//-0.638457 
								   16'b0000001010111011,	//0.341071 
								   16'b1111011100101001,	//-1.104752 
								   16'b0000100000001010,	//1.005068 
								   16'b1111100000101010,	//-0.979620 
								   16'b0000000000110001,	//0.023828 
								   16'b0000011001011111,	//0.796307 
								   16'b0000110010000010,	//1.563613 
								   16'b0000111010110011,	//1.837166 
								   16'b0000000110000011,	//0.188862 
								   16'b1111010001110000,	//-1.445502 
								   16'b1111010011000111,	//-1.402824 
								   16'b1111100000111110,	//-0.969967 
								   16'b0000101011100111,	//1.362869 
								   16'b1111100000100011,	//-0.982871 
								   16'b0000101000001111,	//1.257139 
								   16'b1111011111001011,	//-1.025900 
								   16'b0000110110111101,	//1.717054 
								   16'b1111101100110011,	//-0.600065 
								   16'b1111011001001011,	//-1.213619 
								   16'b1111100000001001,	//-0.995665 
								   16'b0000001110110111,	//0.464179 
								   16'b1111111100100101,	//-0.106845 
								   16'b1111101101000001,	//-0.593362 
								   16'b0000101010010110,	//1.323315 
								   16'b0000001010111010,	//0.341056 
								   16'b0000000110010111,	//0.198894 
								   16'b0000110101011010,	//1.668775 
								   16'b1111100100100110,	//-0.856644 
								   16'b0000100000111011,	//1.028801 
								   16'b0000100000011111,	//1.014916 
								   16'b1111110000101101,	//-0.478217 
								   16'b0000001000101100,	//0.271287 
								   16'b1111001001101101,	//-1.696583 
								   16'b1111000110111010,	//-1.784200 
								   16'b0000000011111100,	//0.123190 
								   16'b0000100011101111,	//1.116669 
								   16'b0000110111100011,	//1.736043 
								   16'b1111010000101000,	//-1.480375 
								   16'b0000001000110100,	//0.275295 
								   16'b1111111100000101,	//-0.122437 
								   16'b1111000001100010,	//-1.952392 
								   16'b1111101011001010,	//-0.651509 
								   16'b1111010100110001,	//-1.351271 
								   16'b0000100101101011,	//1.177138 
								   16'b1111100111110101,	//-0.755140 
								   16'b0000000011101010,	//0.114133 
								   16'b1111010101001101,	//-1.337405 
								   16'b0000001101000011,	//0.407928 
								   16'b1111100001101010,	//-0.948115 
								   16'b0000010011101110,	//0.616316 
								   16'b0000011000001110,	//0.756858 
								   16'b0000011111110001,	//0.992606 
								   16'b1111111001101011,	//-0.197834 
								   16'b1111001010101111,	//-1.664714 
								   16'b1111011101010100,	//-1.084092 
								   16'b0000110100111010,	//1.653349 
								   16'b1111010011100000,	//-1.390488 
								   16'b0000101001101101,	//1.303268 
								   16'b0000000100111010,	//0.153370 
								   16'b0000111111100000,	//1.984539 
								   16'b1111001010000000,	//-1.687298 
								   16'b1111111000101010,	//-0.229287 
								   16'b1111001101101010,	//-1.573389 
								   16'b0000111011001000,	//1.847592 
								   16'b1111000000100110,	//-1.981463 
								   16'b0000100011001100,	//1.099642 
								   16'b0000101000100111,	//1.269213 
								   16'b0000101111001100,	//1.474779 
								   16'b1111001010110100,	//-1.662257 
								   16'b1111110011001011,	//-0.400869 
								   16'b1111100001010001,	//-0.960518 
								   16'b0000100110011010,	//1.200274 
								   16'b1111110111001110,	//-0.274345 
								   16'b0000110100100100,	//1.642590 
								   16'b1111010111010010,	//-1.272612 
								   16'b1111100001110001,	//-0.944788 
								   16'b1111010010101000,	//-1.417844 
								   16'b1111010001011011,	//-1.455726 
								   16'b0000101111010001,	//1.477169 
								   16'b0000001010001101,	//0.318818 
								   16'b0000000110011000,	//0.199441 
								   16'b1111010010100011,	//-1.420181 
								   16'b0000101101001100,	//1.412124 
								   16'b0000001111101000,	//0.488221 
								   16'b1111101100111011,	//-0.596190 
								   16'b0000000001101101,	//0.052998 
								   16'b1111110011011100,	//-0.392768 
								   16'b1111001001101110,	//-1.696133 
								   16'b1111011110101101,	//-1.040335 
								   16'b1111001111110010,	//-1.506724 
								   16'b1111010111100011,	//-1.264369 
								   16'b1111011110101110,	//-1.040190 
								   16'b1111110101011010,	//-0.330932 
								   16'b1111000110010111,	//-1.801382 
								   16'b0000110011100011,	//1.610864 
								   16'b0000111000111100,	//1.779149 
								   16'b1111111110110101,	//-0.036544 
								   16'b1111111110101000,	//-0.042989 
								   16'b1111101011001111,	//-0.649122 
								   16'b0000110011001101,	//1.600215 
								   16'b1111101111010001,	//-0.523013 
								   16'b1111001110001111,	//-1.555189 
								   16'b0000100011111000,	//1.121008 
								   16'b1111110001111001,	//-0.441045 
								   16'b1111011110111100,	//-1.033235 
								   16'b1111110011101101,	//-0.384351 
								   16'b1111001100010110,	//-1.614182 
								   16'b1111010000111001,	//-1.472107 
								   16'b0000111000100101,	//1.768202 
								   16'b0000111010011001,	//1.824538 
								   16'b0000001001101000,	//0.300834 
								   16'b1111000111101010,	//-1.760882 
								   16'b1111011110000011,	//-1.060880 
								   16'b1111101101001101,	//-0.587366 
								   16'b0000101001000111,	//1.284776 
								   16'b1111000001111110,	//-1.938386 
								   16'b1111000101100000,	//-1.827905 
								   16'b1111010101101000,	//-1.324040 
								   16'b0000010011000110,	//0.596462 
								   16'b0000011101101010,	//0.926890 
								   16'b0000010010111010,	//0.590984 
								   16'b1111111001101110,	//-0.196305 
								   16'b0000000110000001,	//0.188036 
								   16'b1111100101111011,	//-0.814717 
								   16'b0000011111010101,	//0.978771 
								   16'b1111011000001100,	//-1.244180 
								   16'b0000010111111010,	//0.747102 
								   16'b1111010111011111,	//-1.265955 
								   16'b1111101111001011,	//-0.526062 
								   16'b0000010000000101,	//0.502474 
								   16'b0000100011111000,	//1.120910 
								   16'b1111001010011001,	//-1.675497 
								   16'b0000110110111110,	//1.717544 
								   16'b0000100011010011,	//1.102851 
								   16'b1111111110010100,	//-0.052833 
								   16'b1111110111110011,	//-0.256566 
								   16'b1111111001001100,	//-0.212865 
								   16'b1111100111001110,	//-0.774602 
								   16'b0000000001000110,	//0.034035 
								   16'b0000000001011000,	//0.043086 
								   16'b0000101000101010,	//1.270511 
								   16'b0000100101101111,	//1.179326 
								   16'b0000010010011110,	//0.577273 
								   16'b1111110000011110,	//-0.485562 
								   16'b0000100111111000,	//1.246322 
								   16'b0000000100001101,	//0.131302 
								   16'b1111101100111001,	//-0.597092 
								   16'b0000111000001100,	//1.756006 
								   16'b0000110000001000,	//1.503771 
								   16'b0000000110011011,	//0.200625 
								   16'b0000001111101011,	//0.489900 
								   16'b0000001011001001,	//0.348179 
								   16'b1111011010100110,	//-1.169031 
								   16'b1111100110100100,	//-0.795015 
								   16'b1111111100010010,	//-0.116307 
								   16'b1111011101100000,	//-1.078047 
								   16'b0000101100000101,	//1.377235 
								   16'b1111011000111100,	//-1.220943 
								   16'b1111011100111011,	//-1.096313 
								   16'b1111010101110110,	//-1.317168 
								   16'b1111011101001001,	//-1.089343 
								   16'b1111110111110001,	//-0.257205 
								   16'b1111100111110101,	//-0.755591 
								   16'b0000110110001100,	//1.693519 
								   16'b1111110111000100,	//-0.279170 
								   16'b1111010111101010,	//-1.260735 
								   16'b0000110011110101,	//1.619524 
								   16'b0000111101011010,	//1.918994 
								   16'b1111111000001011,	//-0.244520 
								   16'b1111001110001110,	//-1.555523 
								   16'b1111100001000010,	//-0.967741 
								   16'b1111110100010100,	//-0.365121 
								   16'b0000001100001001,	//0.379584 
								   16'b1111100001100100,	//-0.951153 
								   16'b0000001101001010,	//0.411372 
								   16'b0000011011000010,	//0.844863 
								   16'b1111011100011001,	//-1.113013 
								   16'b1111001111000010,	//-1.530329 
								   16'b1111100101111110,	//-0.813297 
								   16'b1111101000110011,	//-0.724887 
								   16'b1111110110010011,	//-0.303333 
								   16'b0000000001000000,	//0.031433 
								   16'b1111001010111101,	//-1.657937 
								   16'b1111100001100110,	//-0.950071 
								   16'b0000100110100010,	//1.204058 
								   16'b1111000011101111,	//-1.883119 
								   16'b0000110110111001,	//1.715417 
								   16'b0000011101011111,	//0.921323 
								   16'b1111111110100011,	//-0.045564 
								   16'b0000001010000011,	//0.314100 
								   16'b1111011110011000,	//-1.050866 
								   16'b1111111010101111,	//-0.164605 
								   16'b0000111011010010,	//1.852354 
								   16'b0000000101111111,	//0.187223 
								   16'b0000000010101101,	//0.084543 
								   16'b1111011101101001,	//-1.073622 
								   16'b1111111110100101,	//-0.044409 
								   16'b0000001111111000,	//0.496240 
								   16'b0000010110111011,	//0.716542 
								   16'b1111110010101000,	//-0.417939 
								   16'b1111101111000010,	//-0.530253 
								   16'b0000111110011110,	//1.951928 
								   16'b1111000100110101,	//-1.849045 
								   16'b0000110001010011,	//1.540672 
								   16'b0000110100111010,	//1.653147 
								   16'b0000100101111010,	//1.184735 
								   16'b1111001100101001,	//-1.605151 
								   16'b1111100001100001,	//-0.952515 
								   16'b1111101010111011,	//-0.658573 
								   16'b0000010111000000,	//0.718912 
								   16'b1111010001011111,	//-1.453787 
								   16'b0000011100010100,	//0.884910 
								   16'b1111001101101011,	//-1.572953 
								   16'b0000010011101100,	//0.615029 
								   16'b1111111111010000,	//-0.023304 
								   16'b0000100011101110,	//1.116207 
								   16'b0000011011100010,	//0.860148 
								   16'b0000110011101011,	//1.614882 
								   16'b0000110010000010,	//1.563690 
								   16'b1111101010110001,	//-0.663348 
								   16'b0000011001011100,	//0.794983 
								   16'b1111011001010100,	//-1.208761 
								   16'b1111000011111010,	//-1.877836 
								   16'b0000011111001111,	//0.976297 
								   16'b0000000000000000,	//0.000090 
								   16'b1111111101011100,	//-0.080311 
								   16'b0000110011110011,	//1.618889 
								   16'b0000001110000100,	//0.439467 
								   16'b0000001111000100,	//0.470666 
								   16'b0000101110000001,	//1.437769 
								   16'b0000100111000111,	//1.221958 
								   16'b0000001001110101,	//0.306886 
								   16'b1111010111011011,	//-1.268310 
								   16'b1111011110101110,	//-1.040272 
								   16'b0000110001011110,	//1.546048 
								   16'b1111000011101011,	//-1.885303 
								   16'b1111111110101101,	//-0.040394 
								   16'b1111010101100000,	//-1.328291 
								   16'b0000111101010001,	//1.914723 
								   16'b0000011011001110,	//0.850778 
								   16'b0000000000000100,	//0.001886 
								   16'b1111111100010011,	//-0.115647 
								   16'b1111000111101000,	//-1.761525 
								   16'b0000010111010011,	//0.727888 
								   16'b1111000101011100,	//-1.830275 
								   16'b1111001001001001,	//-1.714218 
								   16'b0000000010110001,	//0.086599 
								   16'b1111001100011000,	//-1.613080 
								   16'b0000101000101110,	//1.272594 
								   16'b0000101000101001,	//1.270188 
								   16'b0000011100011110,	//0.889758 
								   16'b1111010011001100,	//-1.400538 
								   16'b0000010100011011,	//0.638421 
								   16'b0000000010011000,	//0.074380 
								   16'b0000111100100011,	//1.891898 
								   16'b0000010011000101,	//0.595966 
								   16'b0000100110011100,	//1.201322 
								   16'b1111111010000110,	//-0.184809 
								   16'b1111110111010110,	//-0.270434 
								   16'b0000101001101001,	//1.301255 
								   16'b1111001010101100,	//-1.666121 
								   16'b1111010001000011,	//-1.467316 
								   16'b1111010110001100,	//-1.306446 
								   16'b1111110010000011,	//-0.436249 
								   16'b0000101010011011,	//1.325519 
								   16'b0000100110110101,	//1.213458 
								   16'b1111000111101111,	//-1.758115 
								   16'b1111110011000111,	//-0.402969 
								   16'b0000000011011100,	//0.107503 
								   16'b1111110101010110,	//-0.332802 
								   16'b0000010100000101,	//0.627440 
								   16'b0000010000011000,	//0.511893 
								   16'b1111100101011000,	//-0.832064 
								   16'b1111110111010000,	//-0.273395 
								   16'b1111000001111111,	//-1.938051 
								   16'b0000111101111101,	//1.936255 
								   16'b1111010101011001,	//-1.331326 
								   16'b1111001101100110,	//-1.575135 
								   16'b1111101111101011,	//-0.510361 
								   16'b1111011001010111,	//-1.207526 
								   16'b1111111110101100,	//-0.041249 
								   16'b1111101011011101,	//-0.642026 
								   16'b0000111001110100,	//1.806522 
								   16'b0000110101110011,	//1.681328 
								   16'b1111000110110000,	//-1.789292 
								   16'b0000011110011101,	//0.951432 
								   16'b1111100010011101,	//-0.923522 
								   16'b1111110110001000,	//-0.308658 
								   16'b0000000110001000,	//0.191484 
								   16'b0000111000101011,	//1.770948 
								   16'b1111110101011110,	//-0.329024 
								   16'b0000111101110101,	//1.932210 
								   16'b1111100110100110,	//-0.794180 
								   16'b0000011001101111,	//0.804395 
								   16'b0000010101010011,	//0.665355 
								   16'b0000000101000001,	//0.156506 
								   16'b0000011001010111,	//0.792422 
								   16'b0000010101010100,	//0.666112 
								   16'b1111010110110011,	//-1.287470 
								   16'b1111010000011001,	//-1.487942 
								   16'b0000111111111000,	//1.996322 
								   16'b1111010101111010,	//-1.315516 
								   16'b1111000100001011,	//-1.869597 
								   16'b0000000111110101,	//0.244799 
								   16'b0000110000111000,	//1.527466 
								   16'b0000010101101010,	//0.676701 
								   16'b1111011000011000,	//-1.238267 
								   16'b1111101111001110,	//-0.524334 
								   16'b1111111010111110,	//-0.157096 
								   16'b0000111101101010,	//1.926552 
								   16'b1111010100000001,	//-1.374380 
								   16'b0000101101100000,	//1.422091 
								   16'b0000010010100010,	//0.579058 
								   16'b1111110000001010,	//-0.494911 
								   16'b1111011000011100,	//-1.236305 
								   16'b1111110110110100,	//-0.286988 
								   16'b1111111101101101,	//-0.071912 
								   16'b1111001111011100,	//-1.517554 
								   16'b0000001011011101,	//0.358030 
								   16'b1111011100111101,	//-1.095249 
								   16'b1111110001001111,	//-0.461524 
								   16'b0000001010101000,	//0.331946 
								   16'b1111100000001111,	//-0.992776 
								   16'b1111100101001011,	//-0.838237 
								   16'b0000001110111111,	//0.468364 
								   16'b1111100001111101,	//-0.938876 
								   16'b0000101001100001,	//1.297505 
								   16'b0000111101110010,	//1.930654 
								   16'b0000011101011110,	//0.920995 
								   16'b1111101100000001,	//-0.624492 
								   16'b0000001010110001,	//0.336277 
								   16'b1111001101110011,	//-1.568924 
								   16'b0000110100000000,	//1.625233 
								   16'b0000110000100110,	//1.518615 
								   16'b0000101000101011,	//1.271042 
								   16'b1111100001011000,	//-0.957088 
								   16'b0000001100000101,	//0.377425 
								   16'b1111000010111000,	//-1.909950 
								   16'b1111110110011100,	//-0.298963 
								   16'b1111101000000010,	//-0.749124 
								   16'b1111010100101011,	//-1.354061 
								   16'b1111010110111000,	//-1.284935 
								   16'b1111110110001000,	//-0.308457 
								   16'b1111001100000100,	//-1.623083 
								   16'b0000001100100111,	//0.394095 
								   16'b1111111100010010,	//-0.116303 
								   16'b0000011001000101,	//0.783797 
								   16'b0000011001100101,	//0.799551 
								   16'b0000010001101111,	//0.554123 
								   16'b1111000100010011,	//-1.865585 
								   16'b1111001000110100,	//-1.724776 
								   16'b1111101000111010,	//-0.721601 
								   16'b0000000011111101,	//0.123457 
								   16'b0000010011110001,	//0.617783 
								   16'b1111110100001011,	//-0.369523 
								   16'b0000101000111101,	//1.279925 
								   16'b0000011011111101,	//0.873436 
								   16'b0000111011111111,	//1.874597 
								   16'b0000000100000001,	//0.125336 
								   16'b1111101001101000,	//-0.699417 
								   16'b1111001101100001,	//-1.577483 
								   16'b0000001110001101,	//0.443835 
								   16'b0000100011101100,	//1.115209 
								   16'b1111110110001101,	//-0.306188 
								   16'b1111001011101000,	//-1.636707 
								   16'b1111100010000111,	//-0.934114 
								   16'b1111010011101011,	//-1.385373 
								   16'b1111100011111110,	//-0.875979 
								   16'b1111111000010101,	//-0.239659 
								   16'b0000000011011110,	//0.108571 
								   16'b1111111010100011,	//-0.170303 
								   16'b0000110000000011,	//1.501486 
								   16'b0000000010010100,	//0.072208 
								   16'b0000111000110010,	//1.774490 
								   16'b0000010001101000,	//0.550836 
								   16'b0000111010100101,	//1.830776 
								   16'b1111011110110100,	//-1.037172 
								   16'b0000010110100011,	//0.704489 
								   16'b1111100101000000,	//-0.843742 
								   16'b0000010101111111,	//0.687233 
								   16'b0000011000111111,	//0.780562 
								   16'b1111001000101101,	//-1.728029 
								   16'b1111100000100111,	//-0.980839 
								   16'b1111011100101011,	//-1.103840 
								   16'b0000010101011111,	//0.671331 
								   16'b0000101100000101,	//1.377569 
								   16'b1111101100000110,	//-0.622150 
								   16'b0000100011111010,	//1.122079 
								   16'b0000010110011100,	//0.701328 
								   16'b1111000000110111,	//-1.973139 
								   16'b0000001101000101,	//0.408682 
								   16'b1111110001100000,	//-0.452915 
								   16'b0000110101010000,	//1.663965 
								   16'b1111000000001001,	//-1.995396 
								   16'b1111111011001100,	//-0.150203 
								   16'b1111110110010100,	//-0.302604 
								   16'b1111111011000000,	//-0.156335 
								   16'b0000100010100101,	//1.080639 
								   16'b1111101001010010,	//-0.710113 
								   16'b0000100100011101,	//1.138957 
								   16'b1111111100010101,	//-0.114571 
								   16'b1111000100100101,	//-1.856949 
								   16'b1111010110100001,	//-1.296502 
								   16'b0000011100011001,	//0.887032 
								   16'b1111111100100111,	//-0.106056 
								   16'b1111010011100011,	//-1.389115 
								   16'b1111101011101010,	//-0.635502 
								   16'b0000001101110000,	//0.429557 
								   16'b1111011000100011,	//-1.233019 
								   16'b0000011110100001,	//0.953707 
								   16'b1111011111000101,	//-1.028602 
								   16'b0000110101011100,	//1.669697 
								   16'b1111100010011100,	//-0.923754 
								   16'b0000100001111111,	//1.062000 
								   16'b1111011000001010,	//-1.245352 
								   16'b1111100100110011,	//-0.850007 
								   16'b1111001011101010,	//-1.635546 
								   16'b0000001001110000,	//0.304838 
								   16'b0000010111011110,	//0.733453 
								   16'b0000000101111110,	//0.186372 
								   16'b1111110110100000,	//-0.297085 
								   16'b0000010010011111,	//0.577771 
								   16'b0000010010111001,	//0.590471 
								   16'b0000010110111011,	//0.716067 
								   16'b0000010001011000,	//0.543147 
								   16'b0000111000111111,	//1.780696 
								   16'b1111011010110000,	//-1.164260 
								   16'b0000011010110010,	//0.837127 
								   16'b1111011110001111,	//-1.055078 
								   16'b1111001111010010,	//-1.522415 
								   16'b0000001101101111,	//0.429216 
								   16'b1111111001101000,	//-0.199449 
								   16'b1111111010101110,	//-0.165098 
								   16'b0000010100101111,	//0.647779 
								   16'b0000100010100110,	//1.081142 
								   16'b1111101100110101,	//-0.599128 
								   16'b0000010100101111,	//0.648038 
								   16'b1111110101010001,	//-0.335366 
								   16'b0000101011110001,	//1.367717 
								   16'b0000101010100111,	//1.331667 
								   16'b1111100000110101,	//-0.974236 
								   16'b0000001110100001,	//0.453843 
								   16'b0000001010100010,	//0.328997 
								   16'b0000000101001110,	//0.162957 
								   16'b0000101111010111,	//1.479764 
								   16'b1111100001111001,	//-0.940884 
								   16'b1111101000101110,	//-0.727704 
								   16'b1111001111010001,	//-1.523142 
								   16'b0000111000010011,	//1.759318 
								   16'b0000010010101000,	//0.582207 
								   16'b1111111101011000,	//-0.082147 
								   16'b0000010001110101,	//0.557268 
								   16'b0000000101101110,	//0.178864 
								   16'b0000010010110111,	//0.589246 
								   16'b0000000101101000,	//0.175544 
								   16'b0000011100010011,	//0.884186 
								   16'b0000000010111000,	//0.089981 
								   16'b0000111111001100,	//1.974818 
								   16'b1111011011111111,	//-1.125293 
								   16'b1111001101100011,	//-1.576807 
								   16'b1111001110000011,	//-1.561210 
								   16'b1111001000001001,	//-1.745635 
								   16'b1111110011110010,	//-0.381680 
								   16'b1111111001011001,	//-0.206508 
								   16'b1111101110110101,	//-0.536735 
								   16'b0000100001101111,	//1.054019 
								   16'b0000010000011000,	//0.511586 
								   16'b0000100010110100,	//1.087922 
								   16'b0000110111011010,	//1.731414 
								   16'b0000111100100001,	//1.890963 
								   16'b1111011000100101,	//-1.231887 
								   16'b1111010001110010,	//-1.444503 
								   16'b0000011001001000,	//0.785065 
								   16'b1111001100000001,	//-1.624720 
								   16'b0000000011010000,	//0.101618 
								   16'b0000000011111001,	//0.121377 
								   16'b0000101110001110,	//1.444559 
								   16'b1111111110000100,	//-0.060587 
								   16'b1111110010010111,	//-0.426175 
								   16'b0000010101111100,	//0.685725 
								   16'b0000011110111000,	//0.965032 
								   16'b0000000010100100,	//0.080210 
								   16'b1111101100100000,	//-0.609149 
								   16'b1111010011001101,	//-1.400011 
								   16'b0000001011000001,	//0.344368 
								   16'b1111100001100011,	//-0.951419 
								   16'b1111000101101100,	//-1.822184 
								   16'b0000100000101000,	//1.019733 
								   16'b1111011111000101,	//-1.028859 
								   16'b1111111000101000,	//-0.230391 
								   16'b0000011000000010,	//0.751184 
								   16'b1111101101111111,	//-0.563087 
								   16'b0000011110010000,	//0.945360 
								   16'b1111110010100001,	//-0.421170 
								   16'b0000010111011111,	//0.733663 
								   16'b0000011010001000,	//0.816190 
								   16'b1111111000100111,	//-0.230778 
								   16'b1111000010100000,	//-1.921690 
								   16'b1111101010010110,	//-0.676568 
								   16'b1111110110010100,	//-0.302762 
								   16'b1111100010100110,	//-0.918918 
								   16'b1111011001001110,	//-1.211785 
								   16'b0000101001001100,	//1.286885 
								   16'b1111110111000010,	//-0.280314 
								   16'b0000110001101001,	//1.551084 
								   16'b1111110010000101,	//-0.435268 
								   16'b0000100010011101,	//1.076458 
								   16'b1111110010110011,	//-0.412834 
								   16'b0000100111011111,	//1.234056 
								   16'b0000100000101010,	//1.020308 
								   16'b1111110000010100,	//-0.490418 
								   16'b1111011011101010,	//-1.135924 
								   16'b0000100101001011,	//1.161629 
								   16'b0000111001100001,	//1.797216 
								   16'b1111101001111011,	//-0.689738 
								   16'b0000010101111011,	//0.685057 
								   16'b1111111000001001,	//-0.245420 
								   16'b0000101010101100,	//1.334002 
								   16'b0000100010011010,	//1.075417 
								   16'b1111010101011010,	//-1.330986 
								   16'b0000101110010101,	//1.447922 
								   16'b0000111110101101,	//1.959489 
								   16'b0000000001110110,	//0.057694 
								   16'b0000110001001100,	//1.537124 
								   16'b0000001011010001,	//0.352104 
								   16'b1111010011110100,	//-1.380991 
								   16'b1111011001100101,	//-1.200549 
								   16'b1111110100000110,	//-0.372181 
								   16'b0000011111110101,	//0.994823 
								   16'b0000101001101011,	//1.302335 
								   16'b0000100101000111,	//1.159852 
								   16'b1111101000110001,	//-0.725903 
								   16'b0000000100010111,	//0.136257 
								   16'b1111001011100001,	//-1.640197 
								   16'b1111001110010011,	//-1.553177 
								   16'b1111010001011101,	//-1.454830 
								   16'b0000010110111000,	//0.714609 
								   16'b1111111111011000,	//-0.019292 
								   16'b1111011000010010,	//-1.241158 
								   16'b1111111111010111,	//-0.019977 
								   16'b1111010010111001,	//-1.409567 
								   16'b1111000111000010,	//-1.780103 
								   16'b0000101100111001,	//1.402851 
								   16'b0000000111110000,	//0.242238 
								   16'b0000110110111111,	//1.718435 
								   16'b0000011001001011,	//0.786669 
								   16'b0000001010100110,	//0.331164 
								   16'b0000101000011000,	//1.261589 
								   16'b0000110000100001,	//1.516056 
								   16'b0000111110100101,	//1.955646 
								   16'b1111000000000100,	//-1.997910 
								   16'b0000101110110010,	//1.461754 
								   16'b0000001110011010,	//0.450266 
								   16'b0000111110101110,	//1.959801 
								   16'b0000000011100011,	//0.110720 
								   16'b1111111101011000,	//-0.081906 
								   16'b0000100110100101,	//1.205390 
								   16'b1111011101001010,	//-1.088628 
								   16'b1111111111110000,	//-0.007623 
								   16'b0000110011010100,	//1.603410 
								   16'b0000001001100100,	//0.298645 
								   16'b0000101100001100,	//1.380713 
								   16'b0000011110100011,	//0.954561 
								   16'b0000001011000000,	//0.343948 
								   16'b1111011111100101,	//-1.013062 
								   16'b0000010101010011,	//0.665665 
								   16'b1111001010101100,	//-1.666069 
								   16'b0000010000001000,	//0.503839 
								   16'b0000010100100110,	//0.643778 
								   16'b0000011101011010,	//0.919007 
								   16'b0000110010000001,	//1.563008 
								   16'b0000111101101111,	//1.929213 
								   16'b0000100010011100,	//1.076116 
								   16'b0000001010011011,	//0.325786 
								   16'b0000110110110101,	//1.713252 
								   16'b0000001010010000,	//0.320361 
								   16'b1111000010001011,	//-1.932068 
								   16'b1111001111011110,	//-1.516562 
								   16'b0000101110011011,	//1.450843 
								   16'b1111111101111111,	//-0.062814 
								   16'b0000101100001001,	//1.379423 
								   16'b1111011010110011,	//-1.162380 
								   16'b0000000110101100,	//0.209165 
								   16'b0000010000101000,	//0.519534 
								   16'b1111000100000110,	//-1.872036 
								   16'b0000001110101100,	//0.458854 
								   16'b1111101110011001,	//-0.550354 
								   16'b1111000110010110,	//-1.801870 
								   16'b1111111110101011,	//-0.041720 
								   16'b1111011000101001,	//-1.229958 
								   16'b1111001111110000,	//-1.507665 
								   16'b1111011010010011,	//-1.178023 
								   16'b1111010010110000,	//-1.413940 
								   16'b1111011000001101,	//-1.243711 
								   16'b1111000101011101,	//-1.829390 
								   16'b0000010001010100,	//0.540792 
								   16'b1111100100000101,	//-0.872533 
								   16'b0000000100111100,	//0.154387 
								   16'b0000011000111111,	//0.780652 
								   16'b1111111111111001,	//-0.003536 
								   16'b0000000100100101,	//0.143204 
								   16'b1111111000111111,	//-0.219267 
								   16'b1111001111110111,	//-1.504271 
								   16'b1111111110110001,	//-0.038571 
								   16'b0000101101001100,	//1.411993 
								   16'b0000101111110111,	//1.495710 
								   16'b1111100010100110,	//-0.918823 
								   16'b1111011010101100,	//-1.166155 
								   16'b0000001000010100,	//0.259918 
								   16'b0000010001111101,	//0.561247 
								   16'b1111110101011000,	//-0.331884 
								   16'b1111011010010111,	//-1.176098 
								   16'b0000111001010101,	//1.791732 
								   16'b1111001010100000,	//-1.671715 
								   16'b1111001101100010,	//-1.577162 
								   16'b1111010010001100,	//-1.431836 
								   16'b1111010101010100,	//-1.334158 
								   16'b0000001111011111,	//0.483835 
								   16'b0000001001011100,	//0.294839 
								   16'b1111000110101011,	//-1.791688 
								   16'b0000110111001100,	//1.724806 
								   16'b0000011101010001,	//0.914647 
								   16'b0000011110011100,	//0.951367 
								   16'b1111001000000111,	//-1.746382 
								   16'b0000101110001001,	//1.441762 
								   16'b0000110111100111,	//1.737620 
								   16'b0000111110000000,	//1.937593 
								   16'b0000101101111100,	//1.435755 
								   16'b0000100100100011,	//1.142236 
								   16'b0000000001101110,	//0.053510 
								   16'b1111010110101111,	//-1.289590 
								   16'b1111110011000001,	//-0.405642 
								   16'b1111010001001001,	//-1.464275 
								   16'b1111000011111101,	//-1.876442 
								   16'b0000111000001101,	//1.756567 
								   16'b1111100110100100,	//-0.794776 
								   16'b1111100101110101,	//-0.817865 
								   16'b1111101010100111,	//-0.668255 
								   16'b1111111011110010,	//-0.131727 
								   16'b0000010010111110,	//0.592794 
								   16'b1111000011001111,	//-1.899087 
								   16'b0000101011110011,	//1.368826 
								   16'b0000000111100100,	//0.236130 
								   16'b0000101101010101,	//1.416400 
								   16'b1111101100100010,	//-0.608483 
								   16'b1111111001000110,	//-0.215893 
								   16'b1111000110111100,	//-1.783042 
								   16'b1111010110101011,	//-1.291570 
								   16'b0000010100110110,	//0.651232 
								   16'b1111101010010110,	//-0.676684 
								   16'b0000110011000000,	//1.593945 
								   16'b1111001111001000,	//-1.527379 
								   16'b0000111110100001,	//1.953672 
								   16'b0000000101001000,	//0.159928 
								   16'b0000011010011111,	//0.827670 
								   16'b0000111111111100,	//1.997966 
								   16'b1111100100110110,	//-0.848603 
								   16'b1111110101000100,	//-0.341910 
								   16'b1111111011100000,	//-0.140640 
								   16'b0000100001110010,	//1.055828 
								   16'b0000101000101111,	//1.272816 
								   16'b1111001100110101,	//-1.599114 
								   16'b1111010110110011,	//-1.287532 
								   16'b1111101110000010,	//-0.561460 
								   16'b1111000111010001,	//-1.773181 
								   16'b0000000010110011,	//0.087543 
								   16'b1111101010111111,	//-0.656604 
								   16'b1111010110011111,	//-1.297324 
								   16'b1111011010110000,	//-1.164213 
								   16'b0000110011110111,	//1.620614 
								   16'b0000010110011101,	//0.701565 
								   16'b1111111011111110,	//-0.126127 
								   16'b0000110100110000,	//1.648530 
								   16'b1111001101010100,	//-1.583954 
								   16'b0000011111011100,	//0.982184 
								   16'b0000011110010000,	//0.945070 
								   16'b0000000111111011,	//0.247446 
								   16'b1111010111100101,	//-1.263224 
								   16'b0000001100011100,	//0.388845 
								   16'b1111100110011001,	//-0.800252 
								   16'b1111010001001011,	//-1.463508 
								   16'b1111011011001110,	//-1.149594 
								   16'b0000110010100011,	//1.579767 
								   16'b1111001001001001,	//-1.714189 
								   16'b1111011111000010,	//-1.030054 
								   16'b1111000110111000,	//-1.784982 
								   16'b1111111000100011,	//-0.233112 
								   16'b1111000001101101,	//-1.946867 
								   16'b0000110010110110,	//1.588765 
								   16'b1111011001001011,	//-1.213367 
								   16'b1111001011111101,	//-1.626518 
								   16'b1111100111010110,	//-0.770532 
								   16'b1111111010011000,	//-0.175769 
								   16'b1111001101000001,	//-1.593322 
								   16'b0000111111011010,	//1.981559 
								   16'b1111101010100001,	//-0.671629 
								   16'b1111100110000100,	//-0.810613 
								   16'b1111000111111100,	//-1.751819 
								   16'b1111100110001011,	//-0.807024 
								   16'b1111000101111100,	//-1.814595 
								   16'b0000000000101100,	//0.021713 
								   16'b0000100001011110,	//1.045704 
								   16'b0000010000110010,	//0.524280 
								   16'b1111001011100000,	//-1.640433 
								   16'b1111001010010110,	//-1.676550 
								   16'b0000100011011111,	//1.108962 
								   16'b0000110011110111,	//1.620539 
								   16'b0000000100010101,	//0.135088 
								   16'b1111001101111110,	//-1.563383 
								   16'b0000101001101101,	//1.303235 
								   16'b1111101011010010,	//-0.647609 
								   16'b1111100101101000,	//-0.824108 
								   16'b0000011111100010,	//0.985254 
								   16'b1111000001010101,	//-1.958654 
								   16'b1111000110001101,	//-1.806211 
								   16'b0000010101100000,	//0.671664 
								   16'b0000001101010000,	//0.413872 
								   16'b0000000011010110,	//0.104410 
								   16'b0000011101011010,	//0.918838 
								   16'b0000011010100010,	//0.829014 
								   16'b0000100100000001,	//1.125508 
								   16'b1111100100110111,	//-0.848092 
								   16'b0000011000101001,	//0.770128 
								   16'b0000000111010000,	//0.226679 
								   16'b1111110010110000,	//-0.413917 
								   16'b1111000111111001};	//-1.753637 
