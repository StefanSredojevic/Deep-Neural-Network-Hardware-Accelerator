//This is actually ROM

module sigmoid_lookup (pi_clka,pi_clkb,pi_ena,pi_enb,pi_addra,pi_addrb,po_doa,po_dob);
    input       pi_clka,pi_clkb,pi_ena,pi_enb;
    input [9:0] pi_addra,pi_addrb;
    output[9:0] po_doa,po_dob;
    


// SIGNALS	
//(*rom_style = "block" *) reg[9:0] data;//Ovo za sad nije potrebno, proveri samo da li ce
                                         //alat za sintezu ovo prepoznati kao brom, ako hoce
                                         //onda samo obrisi ovu liniju koda
reg[9:0] rom[1023:0];
(* dont_touch = "true" *) reg[9:0] po_doa,po_dob;

initial begin
rom[0] = 10'b0100000000; 	rom[1] = 10'b0100000100; 	rom[2] = 10'b0100001000; 	rom[3] = 10'b0100001100; 	
rom[4] = 10'b0100010000; 	rom[5] = 10'b0100010100; 	rom[6] = 10'b0100011000; 	rom[7] = 10'b0100011100; 	
rom[8] = 10'b0100100000; 	rom[9] = 10'b0100100100; 	rom[10] = 10'b0100101000; 	rom[11] = 10'b0100101100; 	
rom[12] = 10'b0100101111; 	rom[13] = 10'b0100110011; 	rom[14] = 10'b0100110111; 	rom[15] = 10'b0100111011; 	
rom[16] = 10'b0100111111; 	rom[17] = 10'b0101000010; 	rom[18] = 10'b0101000110; 	rom[19] = 10'b0101001010; 	
rom[20] = 10'b0101001101; 	rom[21] = 10'b0101010001; 	rom[22] = 10'b0101010101; 	rom[23] = 10'b0101011000; 	
rom[24] = 10'b0101011100; 	rom[25] = 10'b0101011111; 	rom[26] = 10'b0101100011; 	rom[27] = 10'b0101100110; 	
rom[28] = 10'b0101101001; 	rom[29] = 10'b0101101101; 	rom[30] = 10'b0101110000; 	rom[31] = 10'b0101110011; 	
rom[32] = 10'b0101110110; 	rom[33] = 10'b0101111001; 	rom[34] = 10'b0101111101; 	rom[35] = 10'b0110000000; 	
rom[36] = 10'b0110000011; 	rom[37] = 10'b0110000101; 	rom[38] = 10'b0110001000; 	rom[39] = 10'b0110001011; 	
rom[40] = 10'b0110001110; 	rom[41] = 10'b0110010001; 	rom[42] = 10'b0110010011; 	rom[43] = 10'b0110010110; 	
rom[44] = 10'b0110011001; 	rom[45] = 10'b0110011011; 	rom[46] = 10'b0110011110; 	rom[47] = 10'b0110100000; 	
rom[48] = 10'b0110100011; 	rom[49] = 10'b0110100101; 	rom[50] = 10'b0110100111; 	rom[51] = 10'b0110101010; 	
rom[52] = 10'b0110101100; 	rom[53] = 10'b0110101110; 	rom[54] = 10'b0110110000; 	rom[55] = 10'b0110110010; 	
rom[56] = 10'b0110110100; 	rom[57] = 10'b0110110110; 	rom[58] = 10'b0110111000; 	rom[59] = 10'b0110111010; 	
rom[60] = 10'b0110111100; 	rom[61] = 10'b0110111110; 	rom[62] = 10'b0111000000; 	rom[63] = 10'b0111000001; 	
rom[64] = 10'b0111000011; 	rom[65] = 10'b0111000101; 	rom[66] = 10'b0111000110; 	rom[67] = 10'b0111001000; 	
rom[68] = 10'b0111001001; 	rom[69] = 10'b0111001011; 	rom[70] = 10'b0111001100; 	rom[71] = 10'b0111001110; 	
rom[72] = 10'b0111001111; 	rom[73] = 10'b0111010001; 	rom[74] = 10'b0111010010; 	rom[75] = 10'b0111010011; 	
rom[76] = 10'b0111010100; 	rom[77] = 10'b0111010110; 	rom[78] = 10'b0111010111; 	rom[79] = 10'b0111011000; 	
rom[80] = 10'b0111011001; 	rom[81] = 10'b0111011010; 	rom[82] = 10'b0111011011; 	rom[83] = 10'b0111011100; 	
rom[84] = 10'b0111011101; 	rom[85] = 10'b0111011110; 	rom[86] = 10'b0111011111; 	rom[87] = 10'b0111100000; 	
rom[88] = 10'b0111100001; 	rom[89] = 10'b0111100010; 	rom[90] = 10'b0111100011; 	rom[91] = 10'b0111100100; 	
rom[92] = 10'b0111100101; 	rom[93] = 10'b0111100101; 	rom[94] = 10'b0111100110; 	rom[95] = 10'b0111100111; 	
rom[96] = 10'b0111101000; 	rom[97] = 10'b0111101000; 	rom[98] = 10'b0111101001; 	rom[99] = 10'b0111101010; 	
rom[100] = 10'b0111101010; 	rom[101] = 10'b0111101011; 	rom[102] = 10'b0111101100; 	rom[103] = 10'b0111101100; 	
rom[104] = 10'b0111101101; 	rom[105] = 10'b0111101101; 	rom[106] = 10'b0111101110; 	rom[107] = 10'b0111101111; 	
rom[108] = 10'b0111101111; 	rom[109] = 10'b0111110000; 	rom[110] = 10'b0111110000; 	rom[111] = 10'b0111110001; 	
rom[112] = 10'b0111110001; 	rom[113] = 10'b0111110001; 	rom[114] = 10'b0111110010; 	rom[115] = 10'b0111110010; 	
rom[116] = 10'b0111110011; 	rom[117] = 10'b0111110011; 	rom[118] = 10'b0111110011; 	rom[119] = 10'b0111110100; 	
rom[120] = 10'b0111110100; 	rom[121] = 10'b0111110101; 	rom[122] = 10'b0111110101; 	rom[123] = 10'b0111110101; 	
rom[124] = 10'b0111110110; 	rom[125] = 10'b0111110110; 	rom[126] = 10'b0111110110; 	rom[127] = 10'b0111110111; 	
rom[128] = 10'b0111110111; 	rom[129] = 10'b0111110111; 	rom[130] = 10'b0111110111; 	rom[131] = 10'b0111111000; 	
rom[132] = 10'b0111111000; 	rom[133] = 10'b0111111000; 	rom[134] = 10'b0111111000; 	rom[135] = 10'b0111111001; 	
rom[136] = 10'b0111111001; 	rom[137] = 10'b0111111001; 	rom[138] = 10'b0111111001; 	rom[139] = 10'b0111111001; 	
rom[140] = 10'b0111111010; 	rom[141] = 10'b0111111010; 	rom[142] = 10'b0111111010; 	rom[143] = 10'b0111111010; 	
rom[144] = 10'b0111111010; 	rom[145] = 10'b0111111011; 	rom[146] = 10'b0111111011; 	rom[147] = 10'b0111111011; 	
rom[148] = 10'b0111111011; 	rom[149] = 10'b0111111011; 	rom[150] = 10'b0111111011; 	rom[151] = 10'b0111111011; 	
rom[152] = 10'b0111111100; 	rom[153] = 10'b0111111100; 	rom[154] = 10'b0111111100; 	rom[155] = 10'b0111111100; 	
rom[156] = 10'b0111111100; 	rom[157] = 10'b0111111100; 	rom[158] = 10'b0111111100; 	rom[159] = 10'b0111111100; 	
rom[160] = 10'b0111111101; 	rom[161] = 10'b0111111101; 	rom[162] = 10'b0111111101; 	rom[163] = 10'b0111111101; 	
rom[164] = 10'b0111111101; 	rom[165] = 10'b0111111101; 	rom[166] = 10'b0111111101; 	rom[167] = 10'b0111111101; 	
rom[168] = 10'b0111111101; 	rom[169] = 10'b0111111101; 	rom[170] = 10'b0111111101; 	rom[171] = 10'b0111111110; 	
rom[172] = 10'b0111111110; 	rom[173] = 10'b0111111110; 	rom[174] = 10'b0111111110; 	rom[175] = 10'b0111111110; 	
rom[176] = 10'b0111111110; 	rom[177] = 10'b0111111110; 	rom[178] = 10'b0111111110; 	rom[179] = 10'b0111111110; 	
rom[180] = 10'b0111111110; 	rom[181] = 10'b0111111110; 	rom[182] = 10'b0111111110; 	rom[183] = 10'b0111111110; 	
rom[184] = 10'b0111111110; 	rom[185] = 10'b0111111110; 	rom[186] = 10'b0111111110; 	rom[187] = 10'b0111111111; 	
rom[188] = 10'b0111111111; 	rom[189] = 10'b0111111111; 	rom[190] = 10'b0111111111; 	rom[191] = 10'b0111111111; 	
rom[192] = 10'b0111111111; 	rom[193] = 10'b0111111111; 	rom[194] = 10'b0111111111; 	rom[195] = 10'b0111111111; 	
rom[196] = 10'b0111111111; 	rom[197] = 10'b0111111111; 	rom[198] = 10'b0111111111; 	rom[199] = 10'b0111111111; 	
rom[200] = 10'b0111111111; 	rom[201] = 10'b0111111111; 	rom[202] = 10'b0111111111; 	rom[203] = 10'b0111111111; 	
rom[204] = 10'b0111111111; 	rom[205] = 10'b0111111111; 	rom[206] = 10'b0111111111; 	rom[207] = 10'b0111111111; 	
rom[208] = 10'b0111111111; 	rom[209] = 10'b0111111111; 	rom[210] = 10'b0111111111; 	rom[211] = 10'b0111111111; 	
rom[212] = 10'b0111111111; 	rom[213] = 10'b0111111111; 	rom[214] = 10'b0111111111; 	rom[215] = 10'b0111111111; 	
rom[216] = 10'b0111111111; 	rom[217] = 10'b0111111111; 	rom[218] = 10'b0111111111; 	rom[219] = 10'b0111111111; 	
rom[220] = 10'b0111111111; 	rom[221] = 10'b0111111111; 	rom[222] = 10'b1000000000; 	rom[223] = 10'b1000000000; 	
rom[224] = 10'b1000000000; 	rom[225] = 10'b1000000000; 	rom[226] = 10'b1000000000; 	rom[227] = 10'b1000000000; 	
rom[228] = 10'b1000000000; 	rom[229] = 10'b1000000000; 	rom[230] = 10'b1000000000; 	rom[231] = 10'b1000000000; 	
rom[232] = 10'b1000000000; 	rom[233] = 10'b1000000000; 	rom[234] = 10'b1000000000; 	rom[235] = 10'b1000000000; 	
rom[236] = 10'b1000000000; 	rom[237] = 10'b1000000000; 	rom[238] = 10'b1000000000; 	rom[239] = 10'b1000000000; 	
rom[240] = 10'b1000000000; 	rom[241] = 10'b1000000000; 	rom[242] = 10'b1000000000; 	rom[243] = 10'b1000000000; 	
rom[244] = 10'b1000000000; 	rom[245] = 10'b1000000000; 	rom[246] = 10'b1000000000; 	rom[247] = 10'b1000000000; 	
rom[248] = 10'b1000000000; 	rom[249] = 10'b1000000000; 	rom[250] = 10'b1000000000; 	rom[251] = 10'b1000000000; 	
rom[252] = 10'b1000000000; 	rom[253] = 10'b1000000000; 	rom[254] = 10'b1000000000; 	rom[255] = 10'b1000000000; 	
rom[256] = 10'b1000000000; 	rom[257] = 10'b1000000000; 	rom[258] = 10'b1000000000; 	rom[259] = 10'b1000000000; 	
rom[260] = 10'b1000000000; 	rom[261] = 10'b1000000000; 	rom[262] = 10'b1000000000; 	rom[263] = 10'b1000000000; 	
rom[264] = 10'b1000000000; 	rom[265] = 10'b1000000000; 	rom[266] = 10'b1000000000; 	rom[267] = 10'b1000000000; 	
rom[268] = 10'b1000000000; 	rom[269] = 10'b1000000000; 	rom[270] = 10'b1000000000; 	rom[271] = 10'b1000000000; 	
rom[272] = 10'b1000000000; 	rom[273] = 10'b1000000000; 	rom[274] = 10'b1000000000; 	rom[275] = 10'b1000000000; 	
rom[276] = 10'b1000000000; 	rom[277] = 10'b1000000000; 	rom[278] = 10'b1000000000; 	rom[279] = 10'b1000000000; 	
rom[280] = 10'b1000000000; 	rom[281] = 10'b1000000000; 	rom[282] = 10'b1000000000; 	rom[283] = 10'b1000000000; 	
rom[284] = 10'b1000000000; 	rom[285] = 10'b1000000000; 	rom[286] = 10'b1000000000; 	rom[287] = 10'b1000000000; 	
rom[288] = 10'b1000000000; 	rom[289] = 10'b1000000000; 	rom[290] = 10'b1000000000; 	rom[291] = 10'b1000000000; 	
rom[292] = 10'b1000000000; 	rom[293] = 10'b1000000000; 	rom[294] = 10'b1000000000; 	rom[295] = 10'b1000000000; 	
rom[296] = 10'b1000000000; 	rom[297] = 10'b1000000000; 	rom[298] = 10'b1000000000; 	rom[299] = 10'b1000000000; 	
rom[300] = 10'b1000000000; 	rom[301] = 10'b1000000000; 	rom[302] = 10'b1000000000; 	rom[303] = 10'b1000000000; 	
rom[304] = 10'b1000000000; 	rom[305] = 10'b1000000000; 	rom[306] = 10'b1000000000; 	rom[307] = 10'b1000000000; 	
rom[308] = 10'b1000000000; 	rom[309] = 10'b1000000000; 	rom[310] = 10'b1000000000; 	rom[311] = 10'b1000000000; 	
rom[312] = 10'b1000000000; 	rom[313] = 10'b1000000000; 	rom[314] = 10'b1000000000; 	rom[315] = 10'b1000000000; 	
rom[316] = 10'b1000000000; 	rom[317] = 10'b1000000000; 	rom[318] = 10'b1000000000; 	rom[319] = 10'b1000000000; 	
rom[320] = 10'b1000000000; 	rom[321] = 10'b1000000000; 	rom[322] = 10'b1000000000; 	rom[323] = 10'b1000000000; 	
rom[324] = 10'b1000000000; 	rom[325] = 10'b1000000000; 	rom[326] = 10'b1000000000; 	rom[327] = 10'b1000000000; 	
rom[328] = 10'b1000000000; 	rom[329] = 10'b1000000000; 	rom[330] = 10'b1000000000; 	rom[331] = 10'b1000000000; 	
rom[332] = 10'b1000000000; 	rom[333] = 10'b1000000000; 	rom[334] = 10'b1000000000; 	rom[335] = 10'b1000000000; 	
rom[336] = 10'b1000000000; 	rom[337] = 10'b1000000000; 	rom[338] = 10'b1000000000; 	rom[339] = 10'b1000000000; 	
rom[340] = 10'b1000000000; 	rom[341] = 10'b1000000000; 	rom[342] = 10'b1000000000; 	rom[343] = 10'b1000000000; 	
rom[344] = 10'b1000000000; 	rom[345] = 10'b1000000000; 	rom[346] = 10'b1000000000; 	rom[347] = 10'b1000000000; 	
rom[348] = 10'b1000000000; 	rom[349] = 10'b1000000000; 	rom[350] = 10'b1000000000; 	rom[351] = 10'b1000000000; 	
rom[352] = 10'b1000000000; 	rom[353] = 10'b1000000000; 	rom[354] = 10'b1000000000; 	rom[355] = 10'b1000000000; 	
rom[356] = 10'b1000000000; 	rom[357] = 10'b1000000000; 	rom[358] = 10'b1000000000; 	rom[359] = 10'b1000000000; 	
rom[360] = 10'b1000000000; 	rom[361] = 10'b1000000000; 	rom[362] = 10'b1000000000; 	rom[363] = 10'b1000000000; 	
rom[364] = 10'b1000000000; 	rom[365] = 10'b1000000000; 	rom[366] = 10'b1000000000; 	rom[367] = 10'b1000000000; 	
rom[368] = 10'b1000000000; 	rom[369] = 10'b1000000000; 	rom[370] = 10'b1000000000; 	rom[371] = 10'b1000000000; 	
rom[372] = 10'b1000000000; 	rom[373] = 10'b1000000000; 	rom[374] = 10'b1000000000; 	rom[375] = 10'b1000000000; 	
rom[376] = 10'b1000000000; 	rom[377] = 10'b1000000000; 	rom[378] = 10'b1000000000; 	rom[379] = 10'b1000000000; 	
rom[380] = 10'b1000000000; 	rom[381] = 10'b1000000000; 	rom[382] = 10'b1000000000; 	rom[383] = 10'b1000000000; 	
rom[384] = 10'b1000000000; 	rom[385] = 10'b1000000000; 	rom[386] = 10'b1000000000; 	rom[387] = 10'b1000000000; 	
rom[388] = 10'b1000000000; 	rom[389] = 10'b1000000000; 	rom[390] = 10'b1000000000; 	rom[391] = 10'b1000000000; 	
rom[392] = 10'b1000000000; 	rom[393] = 10'b1000000000; 	rom[394] = 10'b1000000000; 	rom[395] = 10'b1000000000; 	
rom[396] = 10'b1000000000; 	rom[397] = 10'b1000000000; 	rom[398] = 10'b1000000000; 	rom[399] = 10'b1000000000; 	
rom[400] = 10'b1000000000; 	rom[401] = 10'b1000000000; 	rom[402] = 10'b1000000000; 	rom[403] = 10'b1000000000; 	
rom[404] = 10'b1000000000; 	rom[405] = 10'b1000000000; 	rom[406] = 10'b1000000000; 	rom[407] = 10'b1000000000; 	
rom[408] = 10'b1000000000; 	rom[409] = 10'b1000000000; 	rom[410] = 10'b1000000000; 	rom[411] = 10'b1000000000; 	
rom[412] = 10'b1000000000; 	rom[413] = 10'b1000000000; 	rom[414] = 10'b1000000000; 	rom[415] = 10'b1000000000; 	
rom[416] = 10'b1000000000; 	rom[417] = 10'b1000000000; 	rom[418] = 10'b1000000000; 	rom[419] = 10'b1000000000; 	
rom[420] = 10'b1000000000; 	rom[421] = 10'b1000000000; 	rom[422] = 10'b1000000000; 	rom[423] = 10'b1000000000; 	
rom[424] = 10'b1000000000; 	rom[425] = 10'b1000000000; 	rom[426] = 10'b1000000000; 	rom[427] = 10'b1000000000; 	
rom[428] = 10'b1000000000; 	rom[429] = 10'b1000000000; 	rom[430] = 10'b1000000000; 	rom[431] = 10'b1000000000; 	
rom[432] = 10'b1000000000; 	rom[433] = 10'b1000000000; 	rom[434] = 10'b1000000000; 	rom[435] = 10'b1000000000; 	
rom[436] = 10'b1000000000; 	rom[437] = 10'b1000000000; 	rom[438] = 10'b1000000000; 	rom[439] = 10'b1000000000; 	
rom[440] = 10'b1000000000; 	rom[441] = 10'b1000000000; 	rom[442] = 10'b1000000000; 	rom[443] = 10'b1000000000; 	
rom[444] = 10'b1000000000; 	rom[445] = 10'b1000000000; 	rom[446] = 10'b1000000000; 	rom[447] = 10'b1000000000; 	
rom[448] = 10'b1000000000; 	rom[449] = 10'b1000000000; 	rom[450] = 10'b1000000000; 	rom[451] = 10'b1000000000; 	
rom[452] = 10'b1000000000; 	rom[453] = 10'b1000000000; 	rom[454] = 10'b1000000000; 	rom[455] = 10'b1000000000; 	
rom[456] = 10'b1000000000; 	rom[457] = 10'b1000000000; 	rom[458] = 10'b1000000000; 	rom[459] = 10'b1000000000; 	
rom[460] = 10'b1000000000; 	rom[461] = 10'b1000000000; 	rom[462] = 10'b1000000000; 	rom[463] = 10'b1000000000; 	
rom[464] = 10'b1000000000; 	rom[465] = 10'b1000000000; 	rom[466] = 10'b1000000000; 	rom[467] = 10'b1000000000; 	
rom[468] = 10'b1000000000; 	rom[469] = 10'b1000000000; 	rom[470] = 10'b1000000000; 	rom[471] = 10'b1000000000; 	
rom[472] = 10'b1000000000; 	rom[473] = 10'b1000000000; 	rom[474] = 10'b1000000000; 	rom[475] = 10'b1000000000; 	
rom[476] = 10'b1000000000; 	rom[477] = 10'b1000000000; 	rom[478] = 10'b1000000000; 	rom[479] = 10'b1000000000; 	
rom[480] = 10'b1000000000; 	rom[481] = 10'b1000000000; 	rom[482] = 10'b1000000000; 	rom[483] = 10'b1000000000; 	
rom[484] = 10'b1000000000; 	rom[485] = 10'b1000000000; 	rom[486] = 10'b1000000000; 	rom[487] = 10'b1000000000; 	
rom[488] = 10'b1000000000; 	rom[489] = 10'b1000000000; 	rom[490] = 10'b1000000000; 	rom[491] = 10'b1000000000; 	
rom[492] = 10'b1000000000; 	rom[493] = 10'b1000000000; 	rom[494] = 10'b1000000000; 	rom[495] = 10'b1000000000; 	
rom[496] = 10'b1000000000; 	rom[497] = 10'b1000000000; 	rom[498] = 10'b1000000000; 	rom[499] = 10'b1000000000; 	
rom[500] = 10'b1000000000; 	rom[501] = 10'b1000000000; 	rom[502] = 10'b1000000000; 	rom[503] = 10'b1000000000; 	
rom[504] = 10'b1000000000; 	rom[505] = 10'b1000000000; 	rom[506] = 10'b1000000000; 	rom[507] = 10'b1000000000; 	
rom[508] = 10'b1000000000; 	rom[509] = 10'b1000000000; 	rom[510] = 10'b1000000000; 	rom[511] = 10'b1000000000; 	
rom[512] = 10'b0011111100; 	rom[513] = 10'b0011111000; 	rom[514] = 10'b0011110100; 	rom[515] = 10'b0011110000; 	
rom[516] = 10'b0011101100; 	rom[517] = 10'b0011101000; 	rom[518] = 10'b0011100100; 	rom[519] = 10'b0011100000; 	
rom[520] = 10'b0011011100; 	rom[521] = 10'b0011011000; 	rom[522] = 10'b0011010100; 	rom[523] = 10'b0011010001; 	
rom[524] = 10'b0011001101; 	rom[525] = 10'b0011001001; 	rom[526] = 10'b0011000101; 	rom[527] = 10'b0011000001; 	
rom[528] = 10'b0010111110; 	rom[529] = 10'b0010111010; 	rom[530] = 10'b0010110110; 	rom[531] = 10'b0010110011; 	
rom[532] = 10'b0010101111; 	rom[533] = 10'b0010101011; 	rom[534] = 10'b0010101000; 	rom[535] = 10'b0010100100; 	
rom[536] = 10'b0010100001; 	rom[537] = 10'b0010011101; 	rom[538] = 10'b0010011010; 	rom[539] = 10'b0010010111; 	
rom[540] = 10'b0010010011; 	rom[541] = 10'b0010010000; 	rom[542] = 10'b0010001101; 	rom[543] = 10'b0010001010; 	
rom[544] = 10'b0010000111; 	rom[545] = 10'b0010000011; 	rom[546] = 10'b0010000000; 	rom[547] = 10'b0001111101; 	
rom[548] = 10'b0001111011; 	rom[549] = 10'b0001111000; 	rom[550] = 10'b0001110101; 	rom[551] = 10'b0001110010; 	
rom[552] = 10'b0001101111; 	rom[553] = 10'b0001101101; 	rom[554] = 10'b0001101010; 	rom[555] = 10'b0001100111; 	
rom[556] = 10'b0001100101; 	rom[557] = 10'b0001100010; 	rom[558] = 10'b0001100000; 	rom[559] = 10'b0001011101; 	
rom[560] = 10'b0001011011; 	rom[561] = 10'b0001011001; 	rom[562] = 10'b0001010110; 	rom[563] = 10'b0001010100; 	
rom[564] = 10'b0001010010; 	rom[565] = 10'b0001010000; 	rom[566] = 10'b0001001110; 	rom[567] = 10'b0001001100; 	
rom[568] = 10'b0001001010; 	rom[569] = 10'b0001001000; 	rom[570] = 10'b0001000110; 	rom[571] = 10'b0001000100; 	
rom[572] = 10'b0001000010; 	rom[573] = 10'b0001000000; 	rom[574] = 10'b0000111111; 	rom[575] = 10'b0000111101; 	
rom[576] = 10'b0000111011; 	rom[577] = 10'b0000111010; 	rom[578] = 10'b0000111000; 	rom[579] = 10'b0000110111; 	
rom[580] = 10'b0000110101; 	rom[581] = 10'b0000110100; 	rom[582] = 10'b0000110010; 	rom[583] = 10'b0000110001; 	
rom[584] = 10'b0000101111; 	rom[585] = 10'b0000101110; 	rom[586] = 10'b0000101101; 	rom[587] = 10'b0000101100; 	
rom[588] = 10'b0000101010; 	rom[589] = 10'b0000101001; 	rom[590] = 10'b0000101000; 	rom[591] = 10'b0000100111; 	
rom[592] = 10'b0000100110; 	rom[593] = 10'b0000100101; 	rom[594] = 10'b0000100100; 	rom[595] = 10'b0000100011; 	
rom[596] = 10'b0000100010; 	rom[597] = 10'b0000100001; 	rom[598] = 10'b0000100000; 	rom[599] = 10'b0000011111; 	
rom[600] = 10'b0000011110; 	rom[601] = 10'b0000011101; 	rom[602] = 10'b0000011100; 	rom[603] = 10'b0000011011; 	
rom[604] = 10'b0000011011; 	rom[605] = 10'b0000011010; 	rom[606] = 10'b0000011001; 	rom[607] = 10'b0000011000; 	
rom[608] = 10'b0000011000; 	rom[609] = 10'b0000010111; 	rom[610] = 10'b0000010110; 	rom[611] = 10'b0000010110; 	
rom[612] = 10'b0000010101; 	rom[613] = 10'b0000010100; 	rom[614] = 10'b0000010100; 	rom[615] = 10'b0000010011; 	
rom[616] = 10'b0000010011; 	rom[617] = 10'b0000010010; 	rom[618] = 10'b0000010001; 	rom[619] = 10'b0000010001; 	
rom[620] = 10'b0000010000; 	rom[621] = 10'b0000010000; 	rom[622] = 10'b0000001111; 	rom[623] = 10'b0000001111; 	
rom[624] = 10'b0000001111; 	rom[625] = 10'b0000001110; 	rom[626] = 10'b0000001110; 	rom[627] = 10'b0000001101; 	
rom[628] = 10'b0000001101; 	rom[629] = 10'b0000001101; 	rom[630] = 10'b0000001100; 	rom[631] = 10'b0000001100; 	
rom[632] = 10'b0000001011; 	rom[633] = 10'b0000001011; 	rom[634] = 10'b0000001011; 	rom[635] = 10'b0000001010; 	
rom[636] = 10'b0000001010; 	rom[637] = 10'b0000001010; 	rom[638] = 10'b0000001001; 	rom[639] = 10'b0000001001; 	
rom[640] = 10'b0000001001; 	rom[641] = 10'b0000001001; 	rom[642] = 10'b0000001000; 	rom[643] = 10'b0000001000; 	
rom[644] = 10'b0000001000; 	rom[645] = 10'b0000001000; 	rom[646] = 10'b0000000111; 	rom[647] = 10'b0000000111; 	
rom[648] = 10'b0000000111; 	rom[649] = 10'b0000000111; 	rom[650] = 10'b0000000111; 	rom[651] = 10'b0000000110; 	
rom[652] = 10'b0000000110; 	rom[653] = 10'b0000000110; 	rom[654] = 10'b0000000110; 	rom[655] = 10'b0000000110; 	
rom[656] = 10'b0000000101; 	rom[657] = 10'b0000000101; 	rom[658] = 10'b0000000101; 	rom[659] = 10'b0000000101; 	
rom[660] = 10'b0000000101; 	rom[661] = 10'b0000000101; 	rom[662] = 10'b0000000101; 	rom[663] = 10'b0000000100; 	
rom[664] = 10'b0000000100; 	rom[665] = 10'b0000000100; 	rom[666] = 10'b0000000100; 	rom[667] = 10'b0000000100; 	
rom[668] = 10'b0000000100; 	rom[669] = 10'b0000000100; 	rom[670] = 10'b0000000100; 	rom[671] = 10'b0000000011; 	
rom[672] = 10'b0000000011; 	rom[673] = 10'b0000000011; 	rom[674] = 10'b0000000011; 	rom[675] = 10'b0000000011; 	
rom[676] = 10'b0000000011; 	rom[677] = 10'b0000000011; 	rom[678] = 10'b0000000011; 	rom[679] = 10'b0000000011; 	
rom[680] = 10'b0000000011; 	rom[681] = 10'b0000000011; 	rom[682] = 10'b0000000010; 	rom[683] = 10'b0000000010; 	
rom[684] = 10'b0000000010; 	rom[685] = 10'b0000000010; 	rom[686] = 10'b0000000010; 	rom[687] = 10'b0000000010; 	
rom[688] = 10'b0000000010; 	rom[689] = 10'b0000000010; 	rom[690] = 10'b0000000010; 	rom[691] = 10'b0000000010; 	
rom[692] = 10'b0000000010; 	rom[693] = 10'b0000000010; 	rom[694] = 10'b0000000010; 	rom[695] = 10'b0000000010; 	
rom[696] = 10'b0000000010; 	rom[697] = 10'b0000000010; 	rom[698] = 10'b0000000001; 	rom[699] = 10'b0000000001; 	
rom[700] = 10'b0000000001; 	rom[701] = 10'b0000000001; 	rom[702] = 10'b0000000001; 	rom[703] = 10'b0000000001; 	
rom[704] = 10'b0000000001; 	rom[705] = 10'b0000000001; 	rom[706] = 10'b0000000001; 	rom[707] = 10'b0000000001; 	
rom[708] = 10'b0000000001; 	rom[709] = 10'b0000000001; 	rom[710] = 10'b0000000001; 	rom[711] = 10'b0000000001; 	
rom[712] = 10'b0000000001; 	rom[713] = 10'b0000000001; 	rom[714] = 10'b0000000001; 	rom[715] = 10'b0000000001; 	
rom[716] = 10'b0000000001; 	rom[717] = 10'b0000000001; 	rom[718] = 10'b0000000001; 	rom[719] = 10'b0000000001; 	
rom[720] = 10'b0000000001; 	rom[721] = 10'b0000000001; 	rom[722] = 10'b0000000001; 	rom[723] = 10'b0000000001; 	
rom[724] = 10'b0000000001; 	rom[725] = 10'b0000000001; 	rom[726] = 10'b0000000001; 	rom[727] = 10'b0000000001; 	
rom[728] = 10'b0000000001; 	rom[729] = 10'b0000000001; 	rom[730] = 10'b0000000001; 	rom[731] = 10'b0000000001; 	
rom[732] = 10'b0000000001; 	rom[733] = 10'b0000000000; 	rom[734] = 10'b0000000000; 	rom[735] = 10'b0000000000; 	
rom[736] = 10'b0000000000; 	rom[737] = 10'b0000000000; 	rom[738] = 10'b0000000000; 	rom[739] = 10'b0000000000; 	
rom[740] = 10'b0000000000; 	rom[741] = 10'b0000000000; 	rom[742] = 10'b0000000000; 	rom[743] = 10'b0000000000; 	
rom[744] = 10'b0000000000; 	rom[745] = 10'b0000000000; 	rom[746] = 10'b0000000000; 	rom[747] = 10'b0000000000; 	
rom[748] = 10'b0000000000; 	rom[749] = 10'b0000000000; 	rom[750] = 10'b0000000000; 	rom[751] = 10'b0000000000; 	
rom[752] = 10'b0000000000; 	rom[753] = 10'b0000000000; 	rom[754] = 10'b0000000000; 	rom[755] = 10'b0000000000; 	
rom[756] = 10'b0000000000; 	rom[757] = 10'b0000000000; 	rom[758] = 10'b0000000000; 	rom[759] = 10'b0000000000; 	
rom[760] = 10'b0000000000; 	rom[761] = 10'b0000000000; 	rom[762] = 10'b0000000000; 	rom[763] = 10'b0000000000; 	
rom[764] = 10'b0000000000; 	rom[765] = 10'b0000000000; 	rom[766] = 10'b0000000000; 	rom[767] = 10'b0000000000; 	
rom[768] = 10'b0000000000; 	rom[769] = 10'b0000000000; 	rom[770] = 10'b0000000000; 	rom[771] = 10'b0000000000; 	
rom[772] = 10'b0000000000; 	rom[773] = 10'b0000000000; 	rom[774] = 10'b0000000000; 	rom[775] = 10'b0000000000; 	
rom[776] = 10'b0000000000; 	rom[777] = 10'b0000000000; 	rom[778] = 10'b0000000000; 	rom[779] = 10'b0000000000; 	
rom[780] = 10'b0000000000; 	rom[781] = 10'b0000000000; 	rom[782] = 10'b0000000000; 	rom[783] = 10'b0000000000; 	
rom[784] = 10'b0000000000; 	rom[785] = 10'b0000000000; 	rom[786] = 10'b0000000000; 	rom[787] = 10'b0000000000; 	
rom[788] = 10'b0000000000; 	rom[789] = 10'b0000000000; 	rom[790] = 10'b0000000000; 	rom[791] = 10'b0000000000; 	
rom[792] = 10'b0000000000; 	rom[793] = 10'b0000000000; 	rom[794] = 10'b0000000000; 	rom[795] = 10'b0000000000; 	
rom[796] = 10'b0000000000; 	rom[797] = 10'b0000000000; 	rom[798] = 10'b0000000000; 	rom[799] = 10'b0000000000; 	
rom[800] = 10'b0000000000; 	rom[801] = 10'b0000000000; 	rom[802] = 10'b0000000000; 	rom[803] = 10'b0000000000; 	
rom[804] = 10'b0000000000; 	rom[805] = 10'b0000000000; 	rom[806] = 10'b0000000000; 	rom[807] = 10'b0000000000; 	
rom[808] = 10'b0000000000; 	rom[809] = 10'b0000000000; 	rom[810] = 10'b0000000000; 	rom[811] = 10'b0000000000; 	
rom[812] = 10'b0000000000; 	rom[813] = 10'b0000000000; 	rom[814] = 10'b0000000000; 	rom[815] = 10'b0000000000; 	
rom[816] = 10'b0000000000; 	rom[817] = 10'b0000000000; 	rom[818] = 10'b0000000000; 	rom[819] = 10'b0000000000; 	
rom[820] = 10'b0000000000; 	rom[821] = 10'b0000000000; 	rom[822] = 10'b0000000000; 	rom[823] = 10'b0000000000; 	
rom[824] = 10'b0000000000; 	rom[825] = 10'b0000000000; 	rom[826] = 10'b0000000000; 	rom[827] = 10'b0000000000; 	
rom[828] = 10'b0000000000; 	rom[829] = 10'b0000000000; 	rom[830] = 10'b0000000000; 	rom[831] = 10'b0000000000; 	
rom[832] = 10'b0000000000; 	rom[833] = 10'b0000000000; 	rom[834] = 10'b0000000000; 	rom[835] = 10'b0000000000; 	
rom[836] = 10'b0000000000; 	rom[837] = 10'b0000000000; 	rom[838] = 10'b0000000000; 	rom[839] = 10'b0000000000; 	
rom[840] = 10'b0000000000; 	rom[841] = 10'b0000000000; 	rom[842] = 10'b0000000000; 	rom[843] = 10'b0000000000; 	
rom[844] = 10'b0000000000; 	rom[845] = 10'b0000000000; 	rom[846] = 10'b0000000000; 	rom[847] = 10'b0000000000; 	
rom[848] = 10'b0000000000; 	rom[849] = 10'b0000000000; 	rom[850] = 10'b0000000000; 	rom[851] = 10'b0000000000; 	
rom[852] = 10'b0000000000; 	rom[853] = 10'b0000000000; 	rom[854] = 10'b0000000000; 	rom[855] = 10'b0000000000; 	
rom[856] = 10'b0000000000; 	rom[857] = 10'b0000000000; 	rom[858] = 10'b0000000000; 	rom[859] = 10'b0000000000; 	
rom[860] = 10'b0000000000; 	rom[861] = 10'b0000000000; 	rom[862] = 10'b0000000000; 	rom[863] = 10'b0000000000; 	
rom[864] = 10'b0000000000; 	rom[865] = 10'b0000000000; 	rom[866] = 10'b0000000000; 	rom[867] = 10'b0000000000; 	
rom[868] = 10'b0000000000; 	rom[869] = 10'b0000000000; 	rom[870] = 10'b0000000000; 	rom[871] = 10'b0000000000; 	
rom[872] = 10'b0000000000; 	rom[873] = 10'b0000000000; 	rom[874] = 10'b0000000000; 	rom[875] = 10'b0000000000; 	
rom[876] = 10'b0000000000; 	rom[877] = 10'b0000000000; 	rom[878] = 10'b0000000000; 	rom[879] = 10'b0000000000; 	
rom[880] = 10'b0000000000; 	rom[881] = 10'b0000000000; 	rom[882] = 10'b0000000000; 	rom[883] = 10'b0000000000; 	
rom[884] = 10'b0000000000; 	rom[885] = 10'b0000000000; 	rom[886] = 10'b0000000000; 	rom[887] = 10'b0000000000; 	
rom[888] = 10'b0000000000; 	rom[889] = 10'b0000000000; 	rom[890] = 10'b0000000000; 	rom[891] = 10'b0000000000; 	
rom[892] = 10'b0000000000; 	rom[893] = 10'b0000000000; 	rom[894] = 10'b0000000000; 	rom[895] = 10'b0000000000; 	
rom[896] = 10'b0000000000; 	rom[897] = 10'b0000000000; 	rom[898] = 10'b0000000000; 	rom[899] = 10'b0000000000; 	
rom[900] = 10'b0000000000; 	rom[901] = 10'b0000000000; 	rom[902] = 10'b0000000000; 	rom[903] = 10'b0000000000; 	
rom[904] = 10'b0000000000; 	rom[905] = 10'b0000000000; 	rom[906] = 10'b0000000000; 	rom[907] = 10'b0000000000; 	
rom[908] = 10'b0000000000; 	rom[909] = 10'b0000000000; 	rom[910] = 10'b0000000000; 	rom[911] = 10'b0000000000; 	
rom[912] = 10'b0000000000; 	rom[913] = 10'b0000000000; 	rom[914] = 10'b0000000000; 	rom[915] = 10'b0000000000; 	
rom[916] = 10'b0000000000; 	rom[917] = 10'b0000000000; 	rom[918] = 10'b0000000000; 	rom[919] = 10'b0000000000; 	
rom[920] = 10'b0000000000; 	rom[921] = 10'b0000000000; 	rom[922] = 10'b0000000000; 	rom[923] = 10'b0000000000; 	
rom[924] = 10'b0000000000; 	rom[925] = 10'b0000000000; 	rom[926] = 10'b0000000000; 	rom[927] = 10'b0000000000; 	
rom[928] = 10'b0000000000; 	rom[929] = 10'b0000000000; 	rom[930] = 10'b0000000000; 	rom[931] = 10'b0000000000; 	
rom[932] = 10'b0000000000; 	rom[933] = 10'b0000000000; 	rom[934] = 10'b0000000000; 	rom[935] = 10'b0000000000; 	
rom[936] = 10'b0000000000; 	rom[937] = 10'b0000000000; 	rom[938] = 10'b0000000000; 	rom[939] = 10'b0000000000; 	
rom[940] = 10'b0000000000; 	rom[941] = 10'b0000000000; 	rom[942] = 10'b0000000000; 	rom[943] = 10'b0000000000; 	
rom[944] = 10'b0000000000; 	rom[945] = 10'b0000000000; 	rom[946] = 10'b0000000000; 	rom[947] = 10'b0000000000; 	
rom[948] = 10'b0000000000; 	rom[949] = 10'b0000000000; 	rom[950] = 10'b0000000000; 	rom[951] = 10'b0000000000; 	
rom[952] = 10'b0000000000; 	rom[953] = 10'b0000000000; 	rom[954] = 10'b0000000000; 	rom[955] = 10'b0000000000; 	
rom[956] = 10'b0000000000; 	rom[957] = 10'b0000000000; 	rom[958] = 10'b0000000000; 	rom[959] = 10'b0000000000; 	
rom[960] = 10'b0000000000; 	rom[961] = 10'b0000000000; 	rom[962] = 10'b0000000000; 	rom[963] = 10'b0000000000; 	
rom[964] = 10'b0000000000; 	rom[965] = 10'b0000000000; 	rom[966] = 10'b0000000000; 	rom[967] = 10'b0000000000; 	
rom[968] = 10'b0000000000; 	rom[969] = 10'b0000000000; 	rom[970] = 10'b0000000000; 	rom[971] = 10'b0000000000; 	
rom[972] = 10'b0000000000; 	rom[973] = 10'b0000000000; 	rom[974] = 10'b0000000000; 	rom[975] = 10'b0000000000; 	
rom[976] = 10'b0000000000; 	rom[977] = 10'b0000000000; 	rom[978] = 10'b0000000000; 	rom[979] = 10'b0000000000; 	
rom[980] = 10'b0000000000; 	rom[981] = 10'b0000000000; 	rom[982] = 10'b0000000000; 	rom[983] = 10'b0000000000; 	
rom[984] = 10'b0000000000; 	rom[985] = 10'b0000000000; 	rom[986] = 10'b0000000000; 	rom[987] = 10'b0000000000; 	
rom[988] = 10'b0000000000; 	rom[989] = 10'b0000000000; 	rom[990] = 10'b0000000000; 	rom[991] = 10'b0000000000; 	
rom[992] = 10'b0000000000; 	rom[993] = 10'b0000000000; 	rom[994] = 10'b0000000000; 	rom[995] = 10'b0000000000; 	
rom[996] = 10'b0000000000; 	rom[997] = 10'b0000000000; 	rom[998] = 10'b0000000000; 	rom[999] = 10'b0000000000; 	
rom[1000] = 10'b0000000000; rom[1001] = 10'b0000000000; rom[1002] = 10'b0000000000; rom[1003] = 10'b0000000000; 	
rom[1004] = 10'b0000000000; rom[1005] = 10'b0000000000; rom[1006] = 10'b0000000000; rom[1007] = 10'b0000000000; 	
rom[1008] = 10'b0000000000; rom[1009] = 10'b0000000000; rom[1010] = 10'b0000000000; rom[1011] = 10'b0000000000; 	
rom[1012] = 10'b0000000000; rom[1013] = 10'b0000000000; rom[1014] = 10'b0000000000; rom[1015] = 10'b0000000000; 	
rom[1016] = 10'b0000000000; rom[1017] = 10'b0000000000; rom[1018] = 10'b0000000000; rom[1019] = 10'b0000000000; 	
rom[1020] = 10'b0000000000; rom[1021] = 10'b0000000000; rom[1022] = 10'b0000000000; rom[1023] = 10'b0000000000;
end

//There is only read option
always @(posedge pi_clka) begin 
	if (pi_ena)
        po_doa <= rom[pi_addra];
end

always @(posedge pi_clkb) begin 
	if (pi_enb)
     	po_dob <= rom[pi_addrb];
end

endmodule : sigmoid_lookup
